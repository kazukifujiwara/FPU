library IEEE;
use IEEE.std_logic_1164.all;

package fsqrt_p is

  component fsqrt is
    port (
      a : in std_logic_vector(31 downto 0);
      s : out std_logic_vector(31 downto 0));
  end component;

end package;


library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_misc.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

library work;
use work.fpu_common_p.all;

entity fsqrt is
  port ( A : in  std_logic_vector(31 downto 0);
         S : out std_logic_vector(31 downto 0));
end entity fsqrt;

architecture blackbox of FSQRT is

  function table(index: std_logic_vector(9 downto 0))
    return std_logic_vector
  is
    variable r : std_logic_vector(63 downto 0);
  begin
    case conv_integer(index) is
      when    0 => r := x"3effe0083f000ffd";
      when    1 => r := x"3effa0383f002ff5";
      when    2 => r := x"3eff60973f004fe5";
      when    3 => r := x"3eff21263f006fcd";
      when    4 => r := x"3efee1e43f008fad";
      when    5 => r := x"3efea2d23f00af86";
      when    6 => r := x"3efe63ed3f00cf56";
      when    7 => r := x"3efe25383f00ef1f";
      when    8 => r := x"3efde6b03f010edf";
      when    9 => r := x"3efda8573f012e98";
      when   10 => r := x"3efd6a2b3f014e4a";
      when   11 => r := x"3efd2c2e3f016df3";
      when   12 => r := x"3efcee5d3f018d95";
      when   13 => r := x"3efcb0ba3f01ad2f";
      when   14 => r := x"3efc73443f01ccc1";
      when   15 => r := x"3efc35fa3f01ec4b";
      when   16 => r := x"3efbf8dd3f020bce";
      when   17 => r := x"3efbbbed3f022b4a";
      when   18 => r := x"3efb7f283f024abd";
      when   19 => r := x"3efb42903f026a29";
      when   20 => r := x"3efb06233f02898e";
      when   21 => r := x"3efac9e13f02a8eb";
      when   22 => r := x"3efa8dcb3f02c840";
      when   23 => r := x"3efa51e03f02e78e";
      when   24 => r := x"3efa16203f0306d5";
      when   25 => r := x"3ef9da8b3f032614";
      when   26 => r := x"3ef99f203f03454c";
      when   27 => r := x"3ef963e03f03647c";
      when   28 => r := x"3ef928c93f0383a5";
      when   29 => r := x"3ef8eddd3f03a2c6";
      when   30 => r := x"3ef8b31a3f03c1e0";
      when   31 => r := x"3ef878813f03e0f3";
      when   32 => r := x"3ef83e113f03fffe";
      when   33 => r := x"3ef803cb3f041f02";
      when   34 => r := x"3ef7c9ad3f043dff";
      when   35 => r := x"3ef78fb83f045cf5";
      when   36 => r := x"3ef755ec3f047be3";
      when   37 => r := x"3ef71c483f049aca";
      when   38 => r := x"3ef6e2cc3f04b9aa";
      when   39 => r := x"3ef6a9783f04d883";
      when   40 => r := x"3ef6704c3f04f755";
      when   41 => r := x"3ef637483f05161f";
      when   42 => r := x"3ef5fe6c3f0534e2";
      when   43 => r := x"3ef5c5b63f05539f";
      when   44 => r := x"3ef58d283f057254";
      when   45 => r := x"3ef554c13f059102";
      when   46 => r := x"3ef51c813f05afa9";
      when   47 => r := x"3ef4e4673f05ce49";
      when   48 => r := x"3ef4ac743f05ece2";
      when   49 => r := x"3ef474a73f060b74";
      when   50 => r := x"3ef43d003f0629ff";
      when   51 => r := x"3ef4057f3f064883";
      when   52 => r := x"3ef3ce233f066701";
      when   53 => r := x"3ef396ee3f068577";
      when   54 => r := x"3ef35fde3f06a3e6";
      when   55 => r := x"3ef328f33f06c24f";
      when   56 => r := x"3ef2f22d3f06e0b1";
      when   57 => r := x"3ef2bb8c3f06ff0c";
      when   58 => r := x"3ef285103f071d60";
      when   59 => r := x"3ef24eb93f073bad";
      when   60 => r := x"3ef218863f0759f3";
      when   61 => r := x"3ef1e2773f077833";
      when   62 => r := x"3ef1ac8d3f07966c";
      when   63 => r := x"3ef176c63f07b49e";
      when   64 => r := x"3ef141243f07d2ca";
      when   65 => r := x"3ef10ba53f07f0ee";
      when   66 => r := x"3ef0d6493f080f0d";
      when   67 => r := x"3ef0a1113f082d24";
      when   68 => r := x"3ef06bfc3f084b35";
      when   69 => r := x"3ef0370a3f08693f";
      when   70 => r := x"3ef0023b3f088743";
      when   71 => r := x"3eefcd8f3f08a540";
      when   72 => r := x"3eef99063f08c336";
      when   73 => r := x"3eef649f3f08e126";
      when   74 => r := x"3eef305a3f08ff0f";
      when   75 => r := x"3eeefc383f091cf2";
      when   76 => r := x"3eeec8373f093ace";
      when   77 => r := x"3eee94593f0958a4";
      when   78 => r := x"3eee609c3f097673";
      when   79 => r := x"3eee2d003f09943c";
      when   80 => r := x"3eedf9873f09b1ff";
      when   81 => r := x"3eedc62e3f09cfbb";
      when   82 => r := x"3eed92f73f09ed70";
      when   83 => r := x"3eed5fe13f0a0b1f";
      when   84 => r := x"3eed2ceb3f0a28c8";
      when   85 => r := x"3eecfa173f0a466b";
      when   86 => r := x"3eecc7633f0a6407";
      when   87 => r := x"3eec94cf3f0a819c";
      when   88 => r := x"3eec625c3f0a9f2c";
      when   89 => r := x"3eec30093f0abcb5";
      when   90 => r := x"3eebfdd63f0ada38";
      when   91 => r := x"3eebcbc43f0af7b5";
      when   92 => r := x"3eeb99d13f0b152b";
      when   93 => r := x"3eeb67fd3f0b329b";
      when   94 => r := x"3eeb36493f0b5005";
      when   95 => r := x"3eeb04b53f0b6d69";
      when   96 => r := x"3eead3403f0b8ac6";
      when   97 => r := x"3eeaa1ea3f0ba81d";
      when   98 => r := x"3eea70b33f0bc56f";
      when   99 => r := x"3eea3f9b3f0be2ba";
      when  100 => r := x"3eea0ea23f0bfffe";
      when  101 => r := x"3ee9ddc83f0c1d3d";
      when  102 => r := x"3ee9ad0c3f0c3a76";
      when  103 => r := x"3ee97c6e3f0c57a9";
      when  104 => r := x"3ee94bef3f0c74d5";
      when  105 => r := x"3ee91b8e3f0c91fc";
      when  106 => r := x"3ee8eb4b3f0caf1c";
      when  107 => r := x"3ee8bb263f0ccc36";
      when  108 => r := x"3ee88b1f3f0ce94b";
      when  109 => r := x"3ee85b353f0d0659";
      when  110 => r := x"3ee82b693f0d2362";
      when  111 => r := x"3ee7fbbb3f0d4064";
      when  112 => r := x"3ee7cc293f0d5d60";
      when  113 => r := x"3ee79cb53f0d7a57";
      when  114 => r := x"3ee76d5e3f0d9748";
      when  115 => r := x"3ee73e253f0db432";
      when  116 => r := x"3ee70f073f0dd117";
      when  117 => r := x"3ee6e0073f0dedf6";
      when  118 => r := x"3ee6b1233f0e0acf";
      when  119 => r := x"3ee6825c3f0e27a2";
      when  120 => r := x"3ee653b23f0e4470";
      when  121 => r := x"3ee625233f0e6137";
      when  122 => r := x"3ee5f6b13f0e7df9";
      when  123 => r := x"3ee5c85b3f0e9ab5";
      when  124 => r := x"3ee59a203f0eb76b";
      when  125 => r := x"3ee56c023f0ed41c";
      when  126 => r := x"3ee53dff3f0ef0c6";
      when  127 => r := x"3ee510183f0f0d6b";
      when  128 => r := x"3ee4e24d3f0f2a0a";
      when  129 => r := x"3ee4b49d3f0f46a4";
      when  130 => r := x"3ee487083f0f6337";
      when  131 => r := x"3ee4598f3f0f7fc5";
      when  132 => r := x"3ee42c303f0f9c4e";
      when  133 => r := x"3ee3feed3f0fb8d1";
      when  134 => r := x"3ee3d1c53f0fd54e";
      when  135 => r := x"3ee3a4b73f0ff1c5";
      when  136 => r := x"3ee377c43f100e37";
      when  137 => r := x"3ee34aeb3f102aa3";
      when  138 => r := x"3ee31e2d3f10470a";
      when  139 => r := x"3ee2f18a3f10636b";
      when  140 => r := x"3ee2c5013f107fc6";
      when  141 => r := x"3ee298913f109c1c";
      when  142 => r := x"3ee26c3c3f10b86c";
      when  143 => r := x"3ee240013f10d4b7";
      when  144 => r := x"3ee213e03f10f0fc";
      when  145 => r := x"3ee1e7d93f110d3c";
      when  146 => r := x"3ee1bbeb3f112976";
      when  147 => r := x"3ee190173f1145ab";
      when  148 => r := x"3ee1645c3f1161da";
      when  149 => r := x"3ee138bb3f117e04";
      when  150 => r := x"3ee10d333f119a28";
      when  151 => r := x"3ee0e1c53f11b647";
      when  152 => r := x"3ee0b66f3f11d261";
      when  153 => r := x"3ee08b323f11ee75";
      when  154 => r := x"3ee0600f3f120a84";
      when  155 => r := x"3ee035043f12268d";
      when  156 => r := x"3ee00a123f124291";
      when  157 => r := x"3edfdf383f125e8f";
      when  158 => r := x"3edfb4773f127a89";
      when  159 => r := x"3edf89cf3f12967d";
      when  160 => r := x"3edf5f3f3f12b26b";
      when  161 => r := x"3edf34c73f12ce54";
      when  162 => r := x"3edf0a673f12ea38";
      when  163 => r := x"3edee0203f130617";
      when  164 => r := x"3edeb5f03f1321f0";
      when  165 => r := x"3ede8bd93f133dc4";
      when  166 => r := x"3ede61d93f135993";
      when  167 => r := x"3ede37f13f13755d";
      when  168 => r := x"3ede0e203f139121";
      when  169 => r := x"3edde4683f13ace0";
      when  170 => r := x"3eddbac63f13c89a";
      when  171 => r := x"3edd913c3f13e44f";
      when  172 => r := x"3edd67ca3f13ffff";
      when  173 => r := x"3edd3e6e3f141ba9";
      when  174 => r := x"3edd152a3f14374e";
      when  175 => r := x"3edcebfd3f1452ee";
      when  176 => r := x"3edcc2e73f146e89";
      when  177 => r := x"3edc99e73f148a1f";
      when  178 => r := x"3edc70ff3f14a5b0";
      when  179 => r := x"3edc482d3f14c13b";
      when  180 => r := x"3edc1f723f14dcc2";
      when  181 => r := x"3edbf6cd3f14f843";
      when  182 => r := x"3edbce3f3f1513c0";
      when  183 => r := x"3edba5c73f152f37";
      when  184 => r := x"3edb7d663f154aa9";
      when  185 => r := x"3edb551b3f156616";
      when  186 => r := x"3edb2ce63f15817e";
      when  187 => r := x"3edb04c73f159ce1";
      when  188 => r := x"3edadcbe3f15b840";
      when  189 => r := x"3edab4cb3f15d399";
      when  190 => r := x"3eda8cee3f15eeed";
      when  191 => r := x"3eda65263f160a3c";
      when  192 => r := x"3eda3d753f162586";
      when  193 => r := x"3eda15d93f1640cb";
      when  194 => r := x"3ed9ee523f165c0b";
      when  195 => r := x"3ed9c6e13f167747";
      when  196 => r := x"3ed99f853f16927d";
      when  197 => r := x"3ed9783f3f16adaf";
      when  198 => r := x"3ed9510e3f16c8db";
      when  199 => r := x"3ed929f23f16e403";
      when  200 => r := x"3ed902eb3f16ff26";
      when  201 => r := x"3ed8dbf93f171a44";
      when  202 => r := x"3ed8b51c3f17355d";
      when  203 => r := x"3ed88e543f175071";
      when  204 => r := x"3ed867a03f176b80";
      when  205 => r := x"3ed841023f17868b";
      when  206 => r := x"3ed81a783f17a191";
      when  207 => r := x"3ed7f4033f17bc92";
      when  208 => r := x"3ed7cda23f17d78e";
      when  209 => r := x"3ed7a7553f17f285";
      when  210 => r := x"3ed7811d3f180d77";
      when  211 => r := x"3ed75af93f182865";
      when  212 => r := x"3ed734ea3f18434e";
      when  213 => r := x"3ed70eef3f185e32";
      when  214 => r := x"3ed6e9073f187912";
      when  215 => r := x"3ed6c3343f1893ed";
      when  216 => r := x"3ed69d753f18aec3";
      when  217 => r := x"3ed677c93f18c994";
      when  218 => r := x"3ed652313f18e461";
      when  219 => r := x"3ed62cad3f18ff29";
      when  220 => r := x"3ed6073d3f1919ec";
      when  221 => r := x"3ed5e1e13f1934aa";
      when  222 => r := x"3ed5bc973f194f64";
      when  223 => r := x"3ed597623f196a1a";
      when  224 => r := x"3ed572403f1984ca";
      when  225 => r := x"3ed54d313f199f76";
      when  226 => r := x"3ed528353f19ba1e";
      when  227 => r := x"3ed5034d3f19d4c0";
      when  228 => r := x"3ed4de773f19ef5e";
      when  229 => r := x"3ed4b9b53f1a09f8";
      when  230 => r := x"3ed495063f1a248d";
      when  231 => r := x"3ed4706a3f1a3f1d";
      when  232 => r := x"3ed44be13f1a59a9";
      when  233 => r := x"3ed4276a3f1a7430";
      when  234 => r := x"3ed403063f1a8eb3";
      when  235 => r := x"3ed3deb53f1aa931";
      when  236 => r := x"3ed3ba773f1ac3aa";
      when  237 => r := x"3ed3964b3f1ade20";
      when  238 => r := x"3ed372323f1af890";
      when  239 => r := x"3ed34e2b3f1b12fc";
      when  240 => r := x"3ed32a363f1b2d64";
      when  241 => r := x"3ed306543f1b47c7";
      when  242 => r := x"3ed2e2843f1b6225";
      when  243 => r := x"3ed2bec73f1b7c7f";
      when  244 => r := x"3ed29b1b3f1b96d5";
      when  245 => r := x"3ed277823f1bb126";
      when  246 => r := x"3ed253fa3f1bcb73";
      when  247 => r := x"3ed230853f1be5bb";
      when  248 => r := x"3ed20d223f1bffff";
      when  249 => r := x"3ed1e9d03f1c1a3e";
      when  250 => r := x"3ed1c6903f1c3479";
      when  251 => r := x"3ed1a3623f1c4eb0";
      when  252 => r := x"3ed180453f1c68e2";
      when  253 => r := x"3ed15d3b3f1c8310";
      when  254 => r := x"3ed13a413f1c9d3a";
      when  255 => r := x"3ed1175a3f1cb75f";
      when  256 => r := x"3ed0f4833f1cd17f";
      when  257 => r := x"3ed0d1be3f1ceb9c";
      when  258 => r := x"3ed0af0b3f1d05b4";
      when  259 => r := x"3ed08c683f1d1fc8";
      when  260 => r := x"3ed069d73f1d39d7";
      when  261 => r := x"3ed047573f1d53e2";
      when  262 => r := x"3ed024e93f1d6de9";
      when  263 => r := x"3ed0028b3f1d87eb";
      when  264 => r := x"3ecfe03e3f1da1e9";
      when  265 => r := x"3ecfbe023f1dbbe3";
      when  266 => r := x"3ecf9bd73f1dd5d9";
      when  267 => r := x"3ecf79bd3f1defca";
      when  268 => r := x"3ecf57b43f1e09b7";
      when  269 => r := x"3ecf35bb3f1e23a0";
      when  270 => r := x"3ecf13d33f1e3d85";
      when  271 => r := x"3ecef1fc3f1e5765";
      when  272 => r := x"3eced0353f1e7141";
      when  273 => r := x"3eceae7f3f1e8b19";
      when  274 => r := x"3ece8cd93f1ea4ed";
      when  275 => r := x"3ece6b443f1ebebc";
      when  276 => r := x"3ece49bf3f1ed888";
      when  277 => r := x"3ece284a3f1ef24f";
      when  278 => r := x"3ece06e63f1f0c12";
      when  279 => r := x"3ecde5923f1f25d1";
      when  280 => r := x"3ecdc44e3f1f3f8b";
      when  281 => r := x"3ecda31a3f1f5942";
      when  282 => r := x"3ecd81f63f1f72f4";
      when  283 => r := x"3ecd60e23f1f8ca2";
      when  284 => r := x"3ecd3fde3f1fa64c";
      when  285 => r := x"3ecd1eea3f1fbff2";
      when  286 => r := x"3eccfe063f1fd994";
      when  287 => r := x"3eccdd323f1ff332";
      when  288 => r := x"3eccbc6d3f200ccb";
      when  289 => r := x"3ecc9bb83f202661";
      when  290 => r := x"3ecc7b133f203ff2";
      when  291 => r := x"3ecc5a7d3f205980";
      when  292 => r := x"3ecc39f73f207309";
      when  293 => r := x"3ecc19813f208c8e";
      when  294 => r := x"3ecbf91a3f20a60f";
      when  295 => r := x"3ecbd8c23f20bf8c";
      when  296 => r := x"3ecbb8793f20d905";
      when  297 => r := x"3ecb98403f20f27a";
      when  298 => r := x"3ecb78173f210beb";
      when  299 => r := x"3ecb57fc3f212558";
      when  300 => r := x"3ecb37f13f213ec1";
      when  301 => r := x"3ecb17f53f215826";
      when  302 => r := x"3ecaf8073f217187";
      when  303 => r := x"3ecad8293f218ae4";
      when  304 => r := x"3ecab85a3f21a43e";
      when  305 => r := x"3eca989a3f21bd93";
      when  306 => r := x"3eca78e93f21d6e4";
      when  307 => r := x"3eca59463f21f031";
      when  308 => r := x"3eca39b33f22097a";
      when  309 => r := x"3eca1a2e3f2222bf";
      when  310 => r := x"3ec9fab83f223c01";
      when  311 => r := x"3ec9db513f22553e";
      when  312 => r := x"3ec9bbf83f226e77";
      when  313 => r := x"3ec99cae3f2287ad";
      when  314 => r := x"3ec97d723f22a0df";
      when  315 => r := x"3ec95e453f22ba0c";
      when  316 => r := x"3ec93f263f22d336";
      when  317 => r := x"3ec920163f22ec5c";
      when  318 => r := x"3ec901143f23057e";
      when  319 => r := x"3ec8e2203f231e9c";
      when  320 => r := x"3ec8c33b3f2337b7";
      when  321 => r := x"3ec8a4643f2350cd";
      when  322 => r := x"3ec8859b3f2369e0";
      when  323 => r := x"3ec866e03f2382ef";
      when  324 => r := x"3ec848333f239bfa";
      when  325 => r := x"3ec829953f23b501";
      when  326 => r := x"3ec80b043f23ce04";
      when  327 => r := x"3ec7ec823f23e703";
      when  328 => r := x"3ec7ce0d3f23ffff";
      when  329 => r := x"3ec7afa63f2418f7";
      when  330 => r := x"3ec7914d3f2431eb";
      when  331 => r := x"3ec773023f244adb";
      when  332 => r := x"3ec754c53f2463c8";
      when  333 => r := x"3ec736963f247cb0";
      when  334 => r := x"3ec718743f249595";
      when  335 => r := x"3ec6fa603f24ae77";
      when  336 => r := x"3ec6dc593f24c754";
      when  337 => r := x"3ec6be603f24e02e";
      when  338 => r := x"3ec6a0753f24f904";
      when  339 => r := x"3ec682973f2511d6";
      when  340 => r := x"3ec664c63f252aa4";
      when  341 => r := x"3ec647033f25436f";
      when  342 => r := x"3ec6294e3f255c36";
      when  343 => r := x"3ec60ba53f2574f9";
      when  344 => r := x"3ec5ee0a3f258db9";
      when  345 => r := x"3ec5d07c3f25a675";
      when  346 => r := x"3ec5b2fc3f25bf2d";
      when  347 => r := x"3ec595883f25d7e2";
      when  348 => r := x"3ec578223f25f092";
      when  349 => r := x"3ec55ac93f260940";
      when  350 => r := x"3ec53d7d3f2621e9";
      when  351 => r := x"3ec5203e3f263a8f";
      when  352 => r := x"3ec5030c3f265331";
      when  353 => r := x"3ec4e5e73f266bd0";
      when  354 => r := x"3ec4c8cf3f26846b";
      when  355 => r := x"3ec4abc43f269d02";
      when  356 => r := x"3ec48ec53f26b596";
      when  357 => r := x"3ec471d43f26ce26";
      when  358 => r := x"3ec454ef3f26e6b2";
      when  359 => r := x"3ec438173f26ff3b";
      when  360 => r := x"3ec41b4b3f2717c0";
      when  361 => r := x"3ec3fe8c3f273042";
      when  362 => r := x"3ec3e1da3f2748c0";
      when  363 => r := x"3ec3c5353f27613a";
      when  364 => r := x"3ec3a89c3f2779b1";
      when  365 => r := x"3ec38c0f3f279224";
      when  366 => r := x"3ec36f8f3f27aa94";
      when  367 => r := x"3ec3531c3f27c300";
      when  368 => r := x"3ec336b53f27db69";
      when  369 => r := x"3ec31a5a3f27f3ce";
      when  370 => r := x"3ec2fe0c3f280c2f";
      when  371 => r := x"3ec2e1ca3f28248d";
      when  372 => r := x"3ec2c5943f283ce8";
      when  373 => r := x"3ec2a96a3f28553f";
      when  374 => r := x"3ec28d4d3f286d92";
      when  375 => r := x"3ec2713c3f2885e2";
      when  376 => r := x"3ec255363f289e2f";
      when  377 => r := x"3ec2393d3f28b677";
      when  378 => r := x"3ec21d513f28cebd";
      when  379 => r := x"3ec201703f28e6ff";
      when  380 => r := x"3ec1e59b3f28ff3d";
      when  381 => r := x"3ec1c9d23f291778";
      when  382 => r := x"3ec1ae153f292fb0";
      when  383 => r := x"3ec192643f2947e4";
      when  384 => r := x"3ec176bf3f296014";
      when  385 => r := x"3ec15b253f297841";
      when  386 => r := x"3ec13f983f29906b";
      when  387 => r := x"3ec124163f29a891";
      when  388 => r := x"3ec108a03f29c0b4";
      when  389 => r := x"3ec0ed353f29d8d3";
      when  390 => r := x"3ec0d1d73f29f0ef";
      when  391 => r := x"3ec0b6833f2a0908";
      when  392 => r := x"3ec09b3c3f2a211d";
      when  393 => r := x"3ec080003f2a392f";
      when  394 => r := x"3ec064d03f2a513d";
      when  395 => r := x"3ec049ab3f2a6948";
      when  396 => r := x"3ec02e913f2a814f";
      when  397 => r := x"3ec013833f2a9954";
      when  398 => r := x"3ebff8813f2ab154";
      when  399 => r := x"3ebfdd8a3f2ac952";
      when  400 => r := x"3ebfc29e3f2ae14c";
      when  401 => r := x"3ebfa7bd3f2af942";
      when  402 => r := x"3ebf8ce83f2b1136";
      when  403 => r := x"3ebf721e3f2b2926";
      when  404 => r := x"3ebf57603f2b4112";
      when  405 => r := x"3ebf3cac3f2b58fb";
      when  406 => r := x"3ebf22043f2b70e1";
      when  407 => r := x"3ebf07673f2b88c4";
      when  408 => r := x"3ebeecd43f2ba0a3";
      when  409 => r := x"3ebed24d3f2bb87f";
      when  410 => r := x"3ebeb7d13f2bd058";
      when  411 => r := x"3ebe9d603f2be82d";
      when  412 => r := x"3ebe82fb3f2bffff";
      when  413 => r := x"3ebe689f3f2c17ce";
      when  414 => r := x"3ebe4e4f3f2c2f99";
      when  415 => r := x"3ebe340a3f2c4761";
      when  416 => r := x"3ebe19d03f2c5f26";
      when  417 => r := x"3ebdffa03f2c76e8";
      when  418 => r := x"3ebde57c3f2c8ea6";
      when  419 => r := x"3ebdcb623f2ca661";
      when  420 => r := x"3ebdb1533f2cbe19";
      when  421 => r := x"3ebd974e3f2cd5ce";
      when  422 => r := x"3ebd7d543f2ced7f";
      when  423 => r := x"3ebd63653f2d052d";
      when  424 => r := x"3ebd49813f2d1cd8";
      when  425 => r := x"3ebd2fa73f2d347f";
      when  426 => r := x"3ebd15d83f2d4c24";
      when  427 => r := x"3ebcfc133f2d63c5";
      when  428 => r := x"3ebce2593f2d7b63";
      when  429 => r := x"3ebcc8a93f2d92fd";
      when  430 => r := x"3ebcaf043f2daa95";
      when  431 => r := x"3ebc95693f2dc229";
      when  432 => r := x"3ebc7bd93f2dd9ba";
      when  433 => r := x"3ebc62533f2df148";
      when  434 => r := x"3ebc48d73f2e08d3";
      when  435 => r := x"3ebc2f663f2e205a";
      when  436 => r := x"3ebc15ff3f2e37df";
      when  437 => r := x"3ebbfca23f2e4f60";
      when  438 => r := x"3ebbe3503f2e66de";
      when  439 => r := x"3ebbca083f2e7e59";
      when  440 => r := x"3ebbb0ca3f2e95d0";
      when  441 => r := x"3ebb97963f2ead45";
      when  442 => r := x"3ebb7e6c3f2ec4b6";
      when  443 => r := x"3ebb654c3f2edc25";
      when  444 => r := x"3ebb4c373f2ef390";
      when  445 => r := x"3ebb332b3f2f0af8";
      when  446 => r := x"3ebb1a2a3f2f225c";
      when  447 => r := x"3ebb01333f2f39be";
      when  448 => r := x"3ebae8453f2f511d";
      when  449 => r := x"3ebacf623f2f6878";
      when  450 => r := x"3ebab6883f2f7fd1";
      when  451 => r := x"3eba9db93f2f9726";
      when  452 => r := x"3eba84f33f2fae78";
      when  453 => r := x"3eba6c373f2fc5c7";
      when  454 => r := x"3eba53853f2fdd13";
      when  455 => r := x"3eba3add3f2ff45c";
      when  456 => r := x"3eba223e3f300ba2";
      when  457 => r := x"3eba09a93f3022e5";
      when  458 => r := x"3eb9f11e3f303a24";
      when  459 => r := x"3eb9d89d3f305161";
      when  460 => r := x"3eb9c0253f30689a";
      when  461 => r := x"3eb9a7b73f307fd1";
      when  462 => r := x"3eb98f533f309704";
      when  463 => r := x"3eb976f83f30ae35";
      when  464 => r := x"3eb95ea73f30c562";
      when  465 => r := x"3eb946603f30dc8c";
      when  466 => r := x"3eb92e213f30f3b4";
      when  467 => r := x"3eb915ed3f310ad8";
      when  468 => r := x"3eb8fdc23f3121f9";
      when  469 => r := x"3eb8e5a03f313917";
      when  470 => r := x"3eb8cd883f315033";
      when  471 => r := x"3eb8b5793f31674b";
      when  472 => r := x"3eb89d743f317e60";
      when  473 => r := x"3eb885783f319572";
      when  474 => r := x"3eb86d853f31ac81";
      when  475 => r := x"3eb8559c3f31c38d";
      when  476 => r := x"3eb83dbc3f31da97";
      when  477 => r := x"3eb825e53f31f19d";
      when  478 => r := x"3eb80e173f3208a0";
      when  479 => r := x"3eb7f6533f321fa0";
      when  480 => r := x"3eb7de983f32369e";
      when  481 => r := x"3eb7c6e63f324d98";
      when  482 => r := x"3eb7af3d3f32648f";
      when  483 => r := x"3eb7979d3f327b84";
      when  484 => r := x"3eb780073f329275";
      when  485 => r := x"3eb768793f32a964";
      when  486 => r := x"3eb750f53f32c04f";
      when  487 => r := x"3eb739793f32d738";
      when  488 => r := x"3eb722073f32ee1e";
      when  489 => r := x"3eb70a9d3f330501";
      when  490 => r := x"3eb6f33d3f331be0";
      when  491 => r := x"3eb6dbe63f3332bd";
      when  492 => r := x"3eb6c4973f334997";
      when  493 => r := x"3eb6ad513f33606f";
      when  494 => r := x"3eb696143f337743";
      when  495 => r := x"3eb67ee13f338e14";
      when  496 => r := x"3eb667b53f33a4e3";
      when  497 => r := x"3eb650933f33bbae";
      when  498 => r := x"3eb6397a3f33d277";
      when  499 => r := x"3eb622693f33e93c";
      when  500 => r := x"3eb60b613f33ffff";
      when  501 => r := x"3eb5f4623f3416bf";
      when  502 => r := x"3eb5dd6b3f342d7c";
      when  503 => r := x"3eb5c67d3f344437";
      when  504 => r := x"3eb5af983f345aee";
      when  505 => r := x"3eb598bc3f3471a3";
      when  506 => r := x"3eb581e83f348854";
      when  507 => r := x"3eb56b1d3f349f03";
      when  508 => r := x"3eb5545a3f34b5af";
      when  509 => r := x"3eb53da03f34cc58";
      when  510 => r := x"3eb526ee3f34e2fe";
      when  511 => r := x"3eb510453f34f9a2";
      when  512 => r := x"3eb4ee583f351b90";
      when  513 => r := x"3eb4c1393f3548c6";
      when  514 => r := x"3eb4943b3f3575f0";
      when  515 => r := x"3eb4675f3f35a310";
      when  516 => r := x"3eb43aa43f35d024";
      when  517 => r := x"3eb40e0b3f35fd2d";
      when  518 => r := x"3eb3e1923f362a2b";
      when  519 => r := x"3eb3b53a3f36571e";
      when  520 => r := x"3eb389033f368406";
      when  521 => r := x"3eb35ced3f36b0e2";
      when  522 => r := x"3eb330f73f36ddb4";
      when  523 => r := x"3eb305213f370a7b";
      when  524 => r := x"3eb2d96c3f373737";
      when  525 => r := x"3eb2add63f3763e8";
      when  526 => r := x"3eb282603f37908e";
      when  527 => r := x"3eb2570a3f37bd29";
      when  528 => r := x"3eb22bd43f37e9b9";
      when  529 => r := x"3eb200bc3f38163f";
      when  530 => r := x"3eb1d5c43f3842ba";
      when  531 => r := x"3eb1aaeb3f386f2a";
      when  532 => r := x"3eb180313f389b8f";
      when  533 => r := x"3eb155963f38c7ea";
      when  534 => r := x"3eb12b193f38f43a";
      when  535 => r := x"3eb100bb3f39207f";
      when  536 => r := x"3eb0d67b3f394cba";
      when  537 => r := x"3eb0ac593f3978eb";
      when  538 => r := x"3eb082553f39a510";
      when  539 => r := x"3eb058703f39d12c";
      when  540 => r := x"3eb02ea83f39fd3d";
      when  541 => r := x"3eb004fd3f3a2943";
      when  542 => r := x"3eafdb713f3a553f";
      when  543 => r := x"3eafb2013f3a8131";
      when  544 => r := x"3eaf88af3f3aad18";
      when  545 => r := x"3eaf5f7a3f3ad8f5";
      when  546 => r := x"3eaf36623f3b04c8";
      when  547 => r := x"3eaf0d663f3b3090";
      when  548 => r := x"3eaee4883f3b5c4f";
      when  549 => r := x"3eaebbc63f3b8803";
      when  550 => r := x"3eae93203f3bb3ad";
      when  551 => r := x"3eae6a973f3bdf4c";
      when  552 => r := x"3eae422a3f3c0ae2";
      when  553 => r := x"3eae19d93f3c366d";
      when  554 => r := x"3eadf1a43f3c61ef";
      when  555 => r := x"3eadc98b3f3c8d66";
      when  556 => r := x"3eada18d3f3cb8d4";
      when  557 => r := x"3ead79ab3f3ce437";
      when  558 => r := x"3ead51e43f3d0f91";
      when  559 => r := x"3ead2a393f3d3ae0";
      when  560 => r := x"3ead02a93f3d6626";
      when  561 => r := x"3eacdb343f3d9161";
      when  562 => r := x"3eacb3da3f3dbc93";
      when  563 => r := x"3eac8c9a3f3de7bb";
      when  564 => r := x"3eac65763f3e12da";
      when  565 => r := x"3eac3e6c3f3e3dee";
      when  566 => r := x"3eac177c3f3e68f9";
      when  567 => r := x"3eabf0a73f3e93fa";
      when  568 => r := x"3eabc9ec3f3ebef1";
      when  569 => r := x"3eaba34c3f3ee9df";
      when  570 => r := x"3eab7cc53f3f14c3";
      when  571 => r := x"3eab56583f3f3f9d";
      when  572 => r := x"3eab30053f3f6a6e";
      when  573 => r := x"3eab09cc3f3f9535";
      when  574 => r := x"3eaae3ac3f3fbff3";
      when  575 => r := x"3eaabda53f3feaa7";
      when  576 => r := x"3eaa97b83f401552";
      when  577 => r := x"3eaa71e53f403ff3";
      when  578 => r := x"3eaa4c2a3f406a8b";
      when  579 => r := x"3eaa26883f409519";
      when  580 => r := x"3eaa00ff3f40bf9e";
      when  581 => r := x"3ea9db8f3f40ea1a";
      when  582 => r := x"3ea9b6383f41148c";
      when  583 => r := x"3ea990f93f413ef5";
      when  584 => r := x"3ea96bd33f416954";
      when  585 => r := x"3ea946c53f4193ab";
      when  586 => r := x"3ea921d03f41bdf8";
      when  587 => r := x"3ea8fcf23f41e83c";
      when  588 => r := x"3ea8d82d3f421276";
      when  589 => r := x"3ea8b3803f423ca8";
      when  590 => r := x"3ea88eea3f4266d0";
      when  591 => r := x"3ea86a6c3f4290ef";
      when  592 => r := x"3ea846063f42bb05";
      when  593 => r := x"3ea821b83f42e512";
      when  594 => r := x"3ea7fd813f430f16";
      when  595 => r := x"3ea7d9613f433911";
      when  596 => r := x"3ea7b5583f436303";
      when  597 => r := x"3ea791673f438cec";
      when  598 => r := x"3ea76d8d3f43b6cc";
      when  599 => r := x"3ea749ca3f43e0a2";
      when  600 => r := x"3ea7261d3f440a70";
      when  601 => r := x"3ea702883f443436";
      when  602 => r := x"3ea6df093f445df2";
      when  603 => r := x"3ea6bba03f4487a5";
      when  604 => r := x"3ea6984f3f44b150";
      when  605 => r := x"3ea675133f44daf1";
      when  606 => r := x"3ea651ee3f45048a";
      when  607 => r := x"3ea62edf3f452e1a";
      when  608 => r := x"3ea60be73f4557a2";
      when  609 => r := x"3ea5e9043f458120";
      when  610 => r := x"3ea5c6373f45aa96";
      when  611 => r := x"3ea5a3803f45d403";
      when  612 => r := x"3ea580df3f45fd68";
      when  613 => r := x"3ea55e543f4626c4";
      when  614 => r := x"3ea53bde3f465017";
      when  615 => r := x"3ea5197e3f467962";
      when  616 => r := x"3ea4f7333f46a2a4";
      when  617 => r := x"3ea4d4fd3f46cbdd";
      when  618 => r := x"3ea4b2dd3f46f50e";
      when  619 => r := x"3ea490d23f471e37";
      when  620 => r := x"3ea46edc3f474757";
      when  621 => r := x"3ea44cfb3f47706e";
      when  622 => r := x"3ea42b2f3f47997d";
      when  623 => r := x"3ea409773f47c284";
      when  624 => r := x"3ea3e7d53f47eb82";
      when  625 => r := x"3ea3c6473f481478";
      when  626 => r := x"3ea3a4cd3f483d65";
      when  627 => r := x"3ea383683f48664a";
      when  628 => r := x"3ea362183f488f27";
      when  629 => r := x"3ea340dc3f48b7fb";
      when  630 => r := x"3ea31fb43f48e0c7";
      when  631 => r := x"3ea2fea03f49098b";
      when  632 => r := x"3ea2dda13f493247";
      when  633 => r := x"3ea2bcb53f495afa";
      when  634 => r := x"3ea29bdd3f4983a5";
      when  635 => r := x"3ea27b1a3f49ac48";
      when  636 => r := x"3ea25a693f49d4e3";
      when  637 => r := x"3ea239cd3f49fd75";
      when  638 => r := x"3ea219443f4a25ff";
      when  639 => r := x"3ea1f8cf3f4a4e82";
      when  640 => r := x"3ea1d86d3f4a76fc";
      when  641 => r := x"3ea1b81f3f4a9f6e";
      when  642 => r := x"3ea197e43f4ac7d8";
      when  643 => r := x"3ea177bc3f4af03a";
      when  644 => r := x"3ea157a83f4b1894";
      when  645 => r := x"3ea137a63f4b40e6";
      when  646 => r := x"3ea117b83f4b6930";
      when  647 => r := x"3ea0f7dc3f4b9172";
      when  648 => r := x"3ea0d8133f4bb9ac";
      when  649 => r := x"3ea0b85e3f4be1de";
      when  650 => r := x"3ea098ba3f4c0a08";
      when  651 => r := x"3ea0792a3f4c322a";
      when  652 => r := x"3ea059ac3f4c5a44";
      when  653 => r := x"3ea03a413f4c8257";
      when  654 => r := x"3ea01ae83f4caa62";
      when  655 => r := x"3e9ffba13f4cd264";
      when  656 => r := x"3e9fdc6d3f4cfa5f";
      when  657 => r := x"3e9fbd4b3f4d2253";
      when  658 => r := x"3e9f9e3b3f4d4a3e";
      when  659 => r := x"3e9f7f3d3f4d7222";
      when  660 => r := x"3e9f60513f4d99fe";
      when  661 => r := x"3e9f41773f4dc1d2";
      when  662 => r := x"3e9f22af3f4de99e";
      when  663 => r := x"3e9f03f93f4e1163";
      when  664 => r := x"3e9ee5553f4e3920";
      when  665 => r := x"3e9ec6c23f4e60d6";
      when  666 => r := x"3e9ea8413f4e8884";
      when  667 => r := x"3e9e89d23f4eb02a";
      when  668 => r := x"3e9e6b743f4ed7c9";
      when  669 => r := x"3e9e4d273f4eff60";
      when  670 => r := x"3e9e2eec3f4f26ef";
      when  671 => r := x"3e9e10c23f4f4e77";
      when  672 => r := x"3e9df2a93f4f75f8";
      when  673 => r := x"3e9dd4a13f4f9d71";
      when  674 => r := x"3e9db6ab3f4fc4e2";
      when  675 => r := x"3e9d98c63f4fec4c";
      when  676 => r := x"3e9d7af13f5013ae";
      when  677 => r := x"3e9d5d2e3f503b09";
      when  678 => r := x"3e9d3f7b3f50625d";
      when  679 => r := x"3e9d21d93f5089a9";
      when  680 => r := x"3e9d04483f50b0ee";
      when  681 => r := x"3e9ce6c83f50d82b";
      when  682 => r := x"3e9cc9583f50ff61";
      when  683 => r := x"3e9cabf83f512690";
      when  684 => r := x"3e9c8eaa3f514db7";
      when  685 => r := x"3e9c716b3f5174d7";
      when  686 => r := x"3e9c543d3f519bf0";
      when  687 => r := x"3e9c371f3f51c302";
      when  688 => r := x"3e9c1a123f51ea0c";
      when  689 => r := x"3e9bfd143f52110f";
      when  690 => r := x"3e9be0273f52380a";
      when  691 => r := x"3e9bc34a3f525eff";
      when  692 => r := x"3e9ba67d3f5285ec";
      when  693 => r := x"3e9b89c03f52acd2";
      when  694 => r := x"3e9b6d133f52d3b1";
      when  695 => r := x"3e9b50753f52fa88";
      when  696 => r := x"3e9b33e83f532159";
      when  697 => r := x"3e9b176a3f534822";
      when  698 => r := x"3e9afafb3f536ee5";
      when  699 => r := x"3e9ade9d3f5395a0";
      when  700 => r := x"3e9ac24e3f53bc54";
      when  701 => r := x"3e9aa60e3f53e301";
      when  702 => r := x"3e9a89de3f5409a7";
      when  703 => r := x"3e9a6dbd3f543046";
      when  704 => r := x"3e9a51ac3f5456de";
      when  705 => r := x"3e9a35aa3f547d6f";
      when  706 => r := x"3e9a19b73f54a3f9";
      when  707 => r := x"3e99fdd33f54ca7c";
      when  708 => r := x"3e99e1fe3f54f0f8";
      when  709 => r := x"3e99c6393f55176d";
      when  710 => r := x"3e99aa823f553ddb";
      when  711 => r := x"3e998edb3f556442";
      when  712 => r := x"3e9973423f558aa2";
      when  713 => r := x"3e9957b83f55b0fc";
      when  714 => r := x"3e993c3d3f55d74e";
      when  715 => r := x"3e9920d13f55fd9a";
      when  716 => r := x"3e9905743f5623df";
      when  717 => r := x"3e98ea253f564a1d";
      when  718 => r := x"3e98cee53f567054";
      when  719 => r := x"3e98b3b33f569684";
      when  720 => r := x"3e9898903f56bcae";
      when  721 => r := x"3e987d7b3f56e2d0";
      when  722 => r := x"3e9862743f5708ec";
      when  723 => r := x"3e98477c3f572f02";
      when  724 => r := x"3e982c933f575510";
      when  725 => r := x"3e9811b73f577b18";
      when  726 => r := x"3e97f6ea3f57a119";
      when  727 => r := x"3e97dc2b3f57c713";
      when  728 => r := x"3e97c17a3f57ed07";
      when  729 => r := x"3e97a6d73f5812f4";
      when  730 => r := x"3e978c423f5838da";
      when  731 => r := x"3e9771bb3f585eba";
      when  732 => r := x"3e9757423f588493";
      when  733 => r := x"3e973cd63f58aa66";
      when  734 => r := x"3e9722793f58d032";
      when  735 => r := x"3e9708293f58f5f7";
      when  736 => r := x"3e96ede83f591bb6";
      when  737 => r := x"3e96d3b33f59416e";
      when  738 => r := x"3e96b98d3f596720";
      when  739 => r := x"3e969f743f598ccb";
      when  740 => r := x"3e9685683f59b26f";
      when  741 => r := x"3e966b6a3f59d80e";
      when  742 => r := x"3e96517a3f59fda5";
      when  743 => r := x"3e9637963f5a2336";
      when  744 => r := x"3e961dc13f5a48c1";
      when  745 => r := x"3e9603f83f5a6e45";
      when  746 => r := x"3e95ea3d3f5a93c3";
      when  747 => r := x"3e95d08f3f5ab93a";
      when  748 => r := x"3e95b6ee3f5adeab";
      when  749 => r := x"3e959d5a3f5b0416";
      when  750 => r := x"3e9583d43f5b297a";
      when  751 => r := x"3e956a5a3f5b4ed8";
      when  752 => r := x"3e9550ee3f5b742f";
      when  753 => r := x"3e95378e3f5b9980";
      when  754 => r := x"3e951e3c3f5bbecb";
      when  755 => r := x"3e9504f63f5be40f";
      when  756 => r := x"3e94ebbd3f5c094d";
      when  757 => r := x"3e94d2913f5c2e85";
      when  758 => r := x"3e94b9713f5c53b7";
      when  759 => r := x"3e94a05f3f5c78e2";
      when  760 => r := x"3e9487583f5c9e07";
      when  761 => r := x"3e946e5f3f5cc326";
      when  762 => r := x"3e9455723f5ce83e";
      when  763 => r := x"3e943c923f5d0d50";
      when  764 => r := x"3e9423be3f5d325c";
      when  765 => r := x"3e940af73f5d5762";
      when  766 => r := x"3e93f23c3f5d7c62";
      when  767 => r := x"3e93d98d3f5da15b";
      when  768 => r := x"3e93c0eb3f5dc64f";
      when  769 => r := x"3e93a8553f5deb3c";
      when  770 => r := x"3e938fcc3f5e1023";
      when  771 => r := x"3e93774e3f5e3504";
      when  772 => r := x"3e935edd3f5e59de";
      when  773 => r := x"3e9346783f5e7eb3";
      when  774 => r := x"3e932e1f3f5ea382";
      when  775 => r := x"3e9315d23f5ec84a";
      when  776 => r := x"3e92fd913f5eed0d";
      when  777 => r := x"3e92e55c3f5f11c9";
      when  778 => r := x"3e92cd333f5f367f";
      when  779 => r := x"3e92b5163f5f5b30";
      when  780 => r := x"3e929d043f5f7fda";
      when  781 => r := x"3e9284ff3f5fa47e";
      when  782 => r := x"3e926d053f5fc91c";
      when  783 => r := x"3e9255183f5fedb5";
      when  784 => r := x"3e923d353f601247";
      when  785 => r := x"3e92255f3f6036d3";
      when  786 => r := x"3e920d943f605b5a";
      when  787 => r := x"3e91f5d53f607fda";
      when  788 => r := x"3e91de213f60a455";
      when  789 => r := x"3e91c6793f60c8c9";
      when  790 => r := x"3e91aedd3f60ed38";
      when  791 => r := x"3e91974b3f6111a1";
      when  792 => r := x"3e917fc63f613603";
      when  793 => r := x"3e91684b3f615a60";
      when  794 => r := x"3e9150dc3f617eb8";
      when  795 => r := x"3e9139793f61a309";
      when  796 => r := x"3e9122203f61c754";
      when  797 => r := x"3e910ad33f61eb9a";
      when  798 => r := x"3e90f3913f620fda";
      when  799 => r := x"3e90dc5a3f623414";
      when  800 => r := x"3e90c52f3f625848";
      when  801 => r := x"3e90ae0e3f627c76";
      when  802 => r := x"3e9096f93f62a09f";
      when  803 => r := x"3e907fee3f62c4c2";
      when  804 => r := x"3e9068ef3f62e8df";
      when  805 => r := x"3e9051fa3f630cf6";
      when  806 => r := x"3e903b113f633108";
      when  807 => r := x"3e9024323f635514";
      when  808 => r := x"3e900d5e3f63791a";
      when  809 => r := x"3e8ff6953f639d1b";
      when  810 => r := x"3e8fdfd73f63c115";
      when  811 => r := x"3e8fc9243f63e50a";
      when  812 => r := x"3e8fb27b3f6408fa";
      when  813 => r := x"3e8f9bdd3f642ce4";
      when  814 => r := x"3e8f854a3f6450c8";
      when  815 => r := x"3e8f6ec13f6474a6";
      when  816 => r := x"3e8f58433f64987f";
      when  817 => r := x"3e8f41d03f64bc53";
      when  818 => r := x"3e8f2b673f64e020";
      when  819 => r := x"3e8f15083f6503e8";
      when  820 => r := x"3e8efeb53f6527ab";
      when  821 => r := x"3e8ee86b3f654b68";
      when  822 => r := x"3e8ed22c3f656f1f";
      when  823 => r := x"3e8ebbf73f6592d1";
      when  824 => r := x"3e8ea5cd3f65b67d";
      when  825 => r := x"3e8e8fad3f65da24";
      when  826 => r := x"3e8e79973f65fdc5";
      when  827 => r := x"3e8e638b3f662160";
      when  828 => r := x"3e8e4d8a3f6644f7";
      when  829 => r := x"3e8e37933f666887";
      when  830 => r := x"3e8e21a63f668c12";
      when  831 => r := x"3e8e0bc33f66af98";
      when  832 => r := x"3e8df5ea3f66d318";
      when  833 => r := x"3e8de01c3f66f693";
      when  834 => r := x"3e8dca573f671a08";
      when  835 => r := x"3e8db49c3f673d78";
      when  836 => r := x"3e8d9eec3f6760e3";
      when  837 => r := x"3e8d89453f678448";
      when  838 => r := x"3e8d73a83f67a7a7";
      when  839 => r := x"3e8d5e153f67cb01";
      when  840 => r := x"3e8d488c3f67ee56";
      when  841 => r := x"3e8d330d3f6811a6";
      when  842 => r := x"3e8d1d983f6834f0";
      when  843 => r := x"3e8d082c3f685835";
      when  844 => r := x"3e8cf2ca3f687b74";
      when  845 => r := x"3e8cdd723f689eae";
      when  846 => r := x"3e8cc8233f68c1e3";
      when  847 => r := x"3e8cb2df3f68e512";
      when  848 => r := x"3e8c9da33f69083c";
      when  849 => r := x"3e8c88723f692b61";
      when  850 => r := x"3e8c734a3f694e80";
      when  851 => r := x"3e8c5e2b3f69719a";
      when  852 => r := x"3e8c49163f6994af";
      when  853 => r := x"3e8c340b3f69b7bf";
      when  854 => r := x"3e8c1f093f69dac9";
      when  855 => r := x"3e8c0a103f69fdcf";
      when  856 => r := x"3e8bf5213f6a20ce";
      when  857 => r := x"3e8be03b3f6a43c9";
      when  858 => r := x"3e8bcb5f3f6a66bf";
      when  859 => r := x"3e8bb68c3f6a89af";
      when  860 => r := x"3e8ba1c23f6aac9a";
      when  861 => r := x"3e8b8d013f6acf80";
      when  862 => r := x"3e8b784a3f6af260";
      when  863 => r := x"3e8b639c3f6b153c";
      when  864 => r := x"3e8b4ef73f6b3812";
      when  865 => r := x"3e8b3a5b3f6b5ae3";
      when  866 => r := x"3e8b25c83f6b7daf";
      when  867 => r := x"3e8b113f3f6ba076";
      when  868 => r := x"3e8afcbe3f6bc338";
      when  869 => r := x"3e8ae8473f6be5f5";
      when  870 => r := x"3e8ad3d93f6c08ac";
      when  871 => r := x"3e8abf733f6c2b5f";
      when  872 => r := x"3e8aab173f6c4e0c";
      when  873 => r := x"3e8a96c33f6c70b4";
      when  874 => r := x"3e8a82793f6c9357";
      when  875 => r := x"3e8a6e373f6cb5f5";
      when  876 => r := x"3e8a59ff3f6cd88e";
      when  877 => r := x"3e8a45cf3f6cfb22";
      when  878 => r := x"3e8a31a83f6d1db1";
      when  879 => r := x"3e8a1d8a3f6d403b";
      when  880 => r := x"3e8a09743f6d62c0";
      when  881 => r := x"3e89f5673f6d8540";
      when  882 => r := x"3e89e1633f6da7bb";
      when  883 => r := x"3e89cd683f6dca31";
      when  884 => r := x"3e89b9763f6deca1";
      when  885 => r := x"3e89a58c3f6e0f0d";
      when  886 => r := x"3e8991aa3f6e3174";
      when  887 => r := x"3e897dd23f6e53d6";
      when  888 => r := x"3e896a013f6e7633";
      when  889 => r := x"3e89563a3f6e988b";
      when  890 => r := x"3e89427b3f6ebade";
      when  891 => r := x"3e892ec43f6edd2c";
      when  892 => r := x"3e891b163f6eff76";
      when  893 => r := x"3e8907713f6f21ba";
      when  894 => r := x"3e88f3d33f6f43f9";
      when  895 => r := x"3e88e03f3f6f6634";
      when  896 => r := x"3e88ccb23f6f886a";
      when  897 => r := x"3e88b92e3f6faa9a";
      when  898 => r := x"3e88a5b33f6fccc6";
      when  899 => r := x"3e88923f3f6feeed";
      when  900 => r := x"3e887ed43f70110f";
      when  901 => r := x"3e886b723f70332d";
      when  902 => r := x"3e8858173f705545";
      when  903 => r := x"3e8844c53f707759";
      when  904 => r := x"3e88317b3f709967";
      when  905 => r := x"3e881e393f70bb71";
      when  906 => r := x"3e880aff3f70dd76";
      when  907 => r := x"3e87f7ce3f70ff77";
      when  908 => r := x"3e87e4a43f712172";
      when  909 => r := x"3e87d1833f714369";
      when  910 => r := x"3e87be693f71655b";
      when  911 => r := x"3e87ab583f718748";
      when  912 => r := x"3e87984f3f71a931";
      when  913 => r := x"3e87854e3f71cb15";
      when  914 => r := x"3e8772543f71ecf3";
      when  915 => r := x"3e875f633f720ece";
      when  916 => r := x"3e874c7a3f7230a3";
      when  917 => r := x"3e8739983f725274";
      when  918 => r := x"3e8726bf3f727440";
      when  919 => r := x"3e8713ed3f729607";
      when  920 => r := x"3e8701233f72b7ca";
      when  921 => r := x"3e86ee613f72d988";
      when  922 => r := x"3e86dba73f72fb41";
      when  923 => r := x"3e86c8f53f731cf6";
      when  924 => r := x"3e86b64a3f733ea6";
      when  925 => r := x"3e86a3a73f736051";
      when  926 => r := x"3e86910c3f7381f7";
      when  927 => r := x"3e867e793f73a399";
      when  928 => r := x"3e866bed3f73c537";
      when  929 => r := x"3e8659693f73e6cf";
      when  930 => r := x"3e8646ec3f740863";
      when  931 => r := x"3e8634783f7429f3";
      when  932 => r := x"3e86220a3f744b7e";
      when  933 => r := x"3e860fa53f746d04";
      when  934 => r := x"3e85fd473f748e85";
      when  935 => r := x"3e85eaf03f74b003";
      when  936 => r := x"3e85d8a13f74d17b";
      when  937 => r := x"3e85c65a3f74f2ef";
      when  938 => r := x"3e85b41a3f75145e";
      when  939 => r := x"3e85a1e13f7535c9";
      when  940 => r := x"3e858fb03f75572f";
      when  941 => r := x"3e857d863f757891";
      when  942 => r := x"3e856b643f7599ee";
      when  943 => r := x"3e8559493f75bb46";
      when  944 => r := x"3e8547353f75dc9b";
      when  945 => r := x"3e8535293f75fdea";
      when  946 => r := x"3e8523243f761f35";
      when  947 => r := x"3e8511273f76407c";
      when  948 => r := x"3e84ff303f7661be";
      when  949 => r := x"3e84ed413f7682fb";
      when  950 => r := x"3e84db5a3f76a434";
      when  951 => r := x"3e84c9793f76c569";
      when  952 => r := x"3e84b7a03f76e699";
      when  953 => r := x"3e84a5cd3f7707c5";
      when  954 => r := x"3e8494023f7728ec";
      when  955 => r := x"3e84823f3f774a0f";
      when  956 => r := x"3e8470823f776b2d";
      when  957 => r := x"3e845ecc3f778c47";
      when  958 => r := x"3e844d1e3f77ad5c";
      when  959 => r := x"3e843b763f77ce6e";
      when  960 => r := x"3e8429d63f77ef7a";
      when  961 => r := x"3e84183d3f781082";
      when  962 => r := x"3e8406aa3f783186";
      when  963 => r := x"3e83f51f3f785286";
      when  964 => r := x"3e83e39b3f787381";
      when  965 => r := x"3e83d21e3f789478";
      when  966 => r := x"3e83c0a73f78b56a";
      when  967 => r := x"3e83af383f78d658";
      when  968 => r := x"3e839dcf3f78f742";
      when  969 => r := x"3e838c6e3f791827";
      when  970 => r := x"3e837b133f793908";
      when  971 => r := x"3e8369bf3f7959e4";
      when  972 => r := x"3e8358723f797abd";
      when  973 => r := x"3e83472c3f799b91";
      when  974 => r := x"3e8335ec3f79bc60";
      when  975 => r := x"3e8324b43f79dd2c";
      when  976 => r := x"3e8313823f79fdf3";
      when  977 => r := x"3e8302573f7a1eb5";
      when  978 => r := x"3e82f1323f7a3f74";
      when  979 => r := x"3e82e0153f7a602e";
      when  980 => r := x"3e82cefe3f7a80e4";
      when  981 => r := x"3e82bdee3f7aa195";
      when  982 => r := x"3e82ace43f7ac243";
      when  983 => r := x"3e829be13f7ae2ec";
      when  984 => r := x"3e828ae53f7b0391";
      when  985 => r := x"3e8279ef3f7b2431";
      when  986 => r := x"3e8269003f7b44ce";
      when  987 => r := x"3e8258183f7b6566";
      when  988 => r := x"3e8247363f7b85fa";
      when  989 => r := x"3e82365a3f7ba689";
      when  990 => r := x"3e8225863f7bc715";
      when  991 => r := x"3e8214b73f7be79c";
      when  992 => r := x"3e8203ef3f7c081f";
      when  993 => r := x"3e81f32e3f7c289e";
      when  994 => r := x"3e81e2733f7c4919";
      when  995 => r := x"3e81d1bf3f7c698f";
      when  996 => r := x"3e81c1113f7c8a02";
      when  997 => r := x"3e81b06a3f7caa70";
      when  998 => r := x"3e819fc83f7ccada";
      when  999 => r := x"3e818f2e3f7ceb40";
      when 1000 => r := x"3e817e993f7d0ba2";
      when 1001 => r := x"3e816e0b3f7d2bff";
      when 1002 => r := x"3e815d843f7d4c59";
      when 1003 => r := x"3e814d023f7d6cae";
      when 1004 => r := x"3e813c873f7d8cff";
      when 1005 => r := x"3e812c133f7dad4c";
      when 1006 => r := x"3e811ba43f7dcd95";
      when 1007 => r := x"3e810b3c3f7dedda";
      when 1008 => r := x"3e80fada3f7e0e1b";
      when 1009 => r := x"3e80ea7f3f7e2e57";
      when 1010 => r := x"3e80da293f7e4e90";
      when 1011 => r := x"3e80c9da3f7e6ec5";
      when 1012 => r := x"3e80b9913f7e8ef5";
      when 1013 => r := x"3e80a94e3f7eaf21";
      when 1014 => r := x"3e8099113f7ecf4a";
      when 1015 => r := x"3e8088db3f7eef6e";
      when 1016 => r := x"3e8078aa3f7f0f8e";
      when 1017 => r := x"3e8068803f7f2faa";
      when 1018 => r := x"3e80585b3f7f4fc2";
      when 1019 => r := x"3e80483d3f7f6fd6";
      when 1020 => r := x"3e8038253f7f8fe6";
      when 1021 => r := x"3e8028133f7faff2";
      when 1022 => r := x"3e8018073f7fcffa";
      when 1023 => r := x"3e8008013f7feffe";
      when others => r := (others => '0');  -- 0 ~ 1023 なのであり得ない。
    end case;
    return r;
  end table;

  component fadd
    port(A : in  std_logic_vector(31 downto 0);
         B : in  std_logic_vector(31 downto 0);
         S : out std_logic_vector(31 downto 0));
  end component;

  component fmul
    port(A : in  std_logic_vector(31 downto 0);
         B : in  std_logic_vector(31 downto 0);
         S : out std_logic_vector(31 downto 0));
  end component;

  constant nan   : std_logic_vector(31 downto 0) := x"7fffffff";
  constant nnan  : std_logic_vector(31 downto 0) := x"ffc00000";
  constant zero  : std_logic_vector(31 downto 0) := x"00000000";
  constant nzero : std_logic_vector(31 downto 0) := x"80000000";
  constant inf   : std_logic_vector(31 downto 0) := x"7f800000";

  signal s1,s2,s3,s4,s5 : std_logic_vector(31 downto 0);

begin

  -- Component Instantiation
  fadd_connect : fadd port map(
    A => s3,
    B => s4,
    S => s5);

  fmul_connect : fmul port map(
    A => s1,
    B => s2,
    S => s3);

  do_fsqrt : process(A, s1, s2, s3, s4, s5)
    variable org      : std_logic_vector(31 downto 0);
    variable result   : std_logic_vector(31 downto 0);
    variable x        : std_logic_vector(31 downto 0);
    variable d        : std_logic_vector(7 downto 0);
    variable index    : std_logic_vector(9 downto 0);
    variable ab_unit  : std_logic_vector(63 downto 0);
    variable ka,kb,temp : std_logic_vector(31 downto 0);   --変更
  begin

    if (is_metavalue(A) or is_metavalue(s3) or is_metavalue(s5)) then
      S <= (others => 'X');
    else
      org := A;

      if org(31) = '1' then
        if org(30 downto 23) = 0 then
          result := nzero;
        else
          result := nnan;
        end if;
      elsif org(30 downto 23) = 0 then
        result := zero;
      elsif org(30 downto 23) = 255 and org(22 downto 0) /= 0 then
        result := nan;
      elsif org = inf then
        result := inf;
      else
        result(31) := '0';
        x := org;
        index := '0' & org(22 downto 14);
        if x(23) = '0' then   -- 指数部のLSBが0のとき(２の奇数乗の場合)
          index(9)  := '1';
          x(30 downto 23) := "10000000";  --128
        else                  -- 指数部のLSBが1のとき(２の偶数乗の場合)
          index(9) := '0';
          x(30 downto 23) := "01111111";  --127
        end if;

        if org(30 downto 23) >= 127 then
          d := org(30 downto 23) - 127;
          d := std_logic_vector(shift_right(unsigned(d), 1));
          result(30 downto 23) := 127 + d;
        else
          d := 127 - org(30 downto 23);
          d := d + 1;
          d := std_logic_vector(shift_right(unsigned(d), 1));
          result(30 downto 23) := 127 - d;
        end if;

        ab_unit := table(index);
        ka := ab_unit(63 downto 32);
        kb := ab_unit(31 downto 0);

        s1 <= ka;
        s2 <= x;
        s4 <= kb;
        temp := s5;

        result(22 downto 0) := temp(22 downto 0);
      end if;

      S <= result;
    end if;
  end process;
end blackbox;

