library ieee;
use ieee.std_logic_1164.all;
use IEEE.numeric_std.all;

library work;
use work.fpu_common_p.all;


package finv_p is

  function finv(a: fpu_data_t) return fpu_data_t;

end package;

package body finv_p is

  type lin is record
    y: unsigned(23 downto 0);
    d: unsigned(23 downto 0);
  end record;

  function finv(a: fpu_data_t)
    return fpu_data_t is

    variable f, g: float_t;
    variable l: lin;
    variable y, d: unsigned(23 downto 0);

  begin

    f := float(a);

    case float_type(a) is
      when NAN =>
        return VAL_NAN;

      when INFORMAL =>
        if f.sign = '0' then
          return VAL_PLUS_INF;
        else
          return VAL_MINUS_INF;
        end if;

      when PLUS_INF =>
        return VAL_PLUS_ZERO;

      when MINUS_INF =>
        return VAL_MINUS_ZERO;

      when PLUS_ZERO =>
        return VAL_PLUS_INF;

      when MINUS_ZERO =>
        return VAL_MINUS_INF;

      when others =>

        l := table(to_integer(f.frac(22 downto 12)));
        g.sign := f.sign;
        g.expt := 253 - g.expt;
        g.frac := resize(l.y + shift_right(l.d * (4096 - f.frac(11 downto 0)), 12), 23);

        return fpu_data(g);
    end case;

  end function;

  type table_t is array(0 to 2047) of lin;

  constant table: table_t := (
    (y => x"ffe003", d => x"001ffd"),
    (y => x"ffc00f", d => x"001ff4"),
    (y => x"ffa023", d => x"001fec"),
    (y => x"ff803f", d => x"001fe4"),
    (y => x"ff6063", d => x"001fdc"),
    (y => x"ff408f", d => x"001fd4"),
    (y => x"ff20c3", d => x"001fcc"),
    (y => x"ff00ff", d => x"001fc4"),
    (y => x"fee142", d => x"001fbd"),
    (y => x"fec18e", d => x"001fb4"),
    (y => x"fea1e1", d => x"001fad"),
    (y => x"fe823c", d => x"001fa5"),
    (y => x"fe629f", d => x"001f9d"),
    (y => x"fe430a", d => x"001f95"),
    (y => x"fe237d", d => x"001f8d"),
    (y => x"fe03f8", d => x"001f85"),
    (y => x"fde47a", d => x"001f7e"),
    (y => x"fdc504", d => x"001f76"),
    (y => x"fda596", d => x"001f6e"),
    (y => x"fd8630", d => x"001f66"),
    (y => x"fd66d2", d => x"001f5e"),
    (y => x"fd477b", d => x"001f57"),
    (y => x"fd282c", d => x"001f4f"),
    (y => x"fd08e5", d => x"001f47"),
    (y => x"fce9a5", d => x"001f40"),
    (y => x"fcca6e", d => x"001f37"),
    (y => x"fcab3e", d => x"001f30"),
    (y => x"fc8c15", d => x"001f29"),
    (y => x"fc6cf5", d => x"001f20"),
    (y => x"fc4ddc", d => x"001f19"),
    (y => x"fc2eca", d => x"001f12"),
    (y => x"fc0fc1", d => x"001f09"),
    (y => x"fbf0be", d => x"001f03"),
    (y => x"fbd1c4", d => x"001efa"),
    (y => x"fbb2d1", d => x"001ef3"),
    (y => x"fb93e6", d => x"001eeb"),
    (y => x"fb7502", d => x"001ee4"),
    (y => x"fb5626", d => x"001edc"),
    (y => x"fb3752", d => x"001ed4"),
    (y => x"fb1885", d => x"001ecd"),
    (y => x"faf9c0", d => x"001ec5"),
    (y => x"fadb02", d => x"001ebe"),
    (y => x"fabc4b", d => x"001eb7"),
    (y => x"fa9d9d", d => x"001eae"),
    (y => x"fa7ef5", d => x"001ea8"),
    (y => x"fa6056", d => x"001e9f"),
    (y => x"fa41bd", d => x"001e99"),
    (y => x"fa232c", d => x"001e91"),
    (y => x"fa04a3", d => x"001e89"),
    (y => x"f9e621", d => x"001e82"),
    (y => x"f9c7a7", d => x"001e7a"),
    (y => x"f9a934", d => x"001e73"),
    (y => x"f98ac8", d => x"001e6c"),
    (y => x"f96c64", d => x"001e64"),
    (y => x"f94e07", d => x"001e5d"),
    (y => x"f92fb2", d => x"001e55"),
    (y => x"f91164", d => x"001e4e"),
    (y => x"f8f31d", d => x"001e47"),
    (y => x"f8d4de", d => x"001e3f"),
    (y => x"f8b6a6", d => x"001e38"),
    (y => x"f89875", d => x"001e31"),
    (y => x"f87a4c", d => x"001e29"),
    (y => x"f85c2a", d => x"001e22"),
    (y => x"f83e0f", d => x"001e1b"),
    (y => x"f81ffc", d => x"001e13"),
    (y => x"f801f0", d => x"001e0c"),
    (y => x"f7e3eb", d => x"001e05"),
    (y => x"f7c5ed", d => x"001dfe"),
    (y => x"f7a7f7", d => x"001df6"),
    (y => x"f78a08", d => x"001def"),
    (y => x"f76c20", d => x"001de8"),
    (y => x"f74e3f", d => x"001de1"),
    (y => x"f73066", d => x"001dd9"),
    (y => x"f71294", d => x"001dd2"),
    (y => x"f6f4c9", d => x"001dcb"),
    (y => x"f6d705", d => x"001dc4"),
    (y => x"f6b948", d => x"001dbd"),
    (y => x"f69b93", d => x"001db5"),
    (y => x"f67de4", d => x"001daf"),
    (y => x"f6603d", d => x"001da7"),
    (y => x"f6429d", d => x"001da0"),
    (y => x"f62504", d => x"001d99"),
    (y => x"f60772", d => x"001d92"),
    (y => x"f5e9e8", d => x"001d8a"),
    (y => x"f5cc64", d => x"001d84"),
    (y => x"f5aee7", d => x"001d7d"),
    (y => x"f59172", d => x"001d75"),
    (y => x"f57403", d => x"001d6f"),
    (y => x"f5569c", d => x"001d67"),
    (y => x"f5393c", d => x"001d60"),
    (y => x"f51be2", d => x"001d5a"),
    (y => x"f4fe90", d => x"001d52"),
    (y => x"f4e145", d => x"001d4b"),
    (y => x"f4c401", d => x"001d44"),
    (y => x"f4a6c3", d => x"001d3e"),
    (y => x"f4898d", d => x"001d36"),
    (y => x"f46c5e", d => x"001d2f"),
    (y => x"f44f35", d => x"001d29"),
    (y => x"f43214", d => x"001d21"),
    (y => x"f414f9", d => x"001d1b"),
    (y => x"f3f7e6", d => x"001d13"),
    (y => x"f3dad9", d => x"001d0d"),
    (y => x"f3bdd4", d => x"001d05"),
    (y => x"f3a0d5", d => x"001cff"),
    (y => x"f383dd", d => x"001cf8"),
    (y => x"f366ec", d => x"001cf1"),
    (y => x"f34a02", d => x"001cea"),
    (y => x"f32d1e", d => x"001ce4"),
    (y => x"f31042", d => x"001cdc"),
    (y => x"f2f36c", d => x"001cd6"),
    (y => x"f2d69e", d => x"001cce"),
    (y => x"f2b9d6", d => x"001cc8"),
    (y => x"f29d15", d => x"001cc1"),
    (y => x"f2805b", d => x"001cba"),
    (y => x"f263a7", d => x"001cb4"),
    (y => x"f246fa", d => x"001cad"),
    (y => x"f22a54", d => x"001ca6"),
    (y => x"f20db5", d => x"001c9f"),
    (y => x"f1f11d", d => x"001c98"),
    (y => x"f1d48b", d => x"001c92"),
    (y => x"f1b801", d => x"001c8a"),
    (y => x"f19b7c", d => x"001c85"),
    (y => x"f17eff", d => x"001c7d"),
    (y => x"f16288", d => x"001c77"),
    (y => x"f14618", d => x"001c70"),
    (y => x"f129af", d => x"001c69"),
    (y => x"f10d4c", d => x"001c63"),
    (y => x"f0f0f1", d => x"001c5b"),
    (y => x"f0d49b", d => x"001c56"),
    (y => x"f0b84d", d => x"001c4e"),
    (y => x"f09c05", d => x"001c48"),
    (y => x"f07fc3", d => x"001c42"),
    (y => x"f06389", d => x"001c3a"),
    (y => x"f04755", d => x"001c34"),
    (y => x"f02b27", d => x"001c2e"),
    (y => x"f00f01", d => x"001c26"),
    (y => x"eff2e0", d => x"001c21"),
    (y => x"efd6c7", d => x"001c19"),
    (y => x"efbab4", d => x"001c13"),
    (y => x"ef9ea7", d => x"001c0d"),
    (y => x"ef82a1", d => x"001c06"),
    (y => x"ef66a2", d => x"001bff"),
    (y => x"ef4aa9", d => x"001bf9"),
    (y => x"ef2eb7", d => x"001bf2"),
    (y => x"ef12cb", d => x"001bec"),
    (y => x"eef6e6", d => x"001be5"),
    (y => x"eedb07", d => x"001bdf"),
    (y => x"eebf2f", d => x"001bd8"),
    (y => x"eea35d", d => x"001bd2"),
    (y => x"ee8792", d => x"001bcb"),
    (y => x"ee6bcd", d => x"001bc5"),
    (y => x"ee500e", d => x"001bbf"),
    (y => x"ee3457", d => x"001bb7"),
    (y => x"ee18a5", d => x"001bb2"),
    (y => x"edfcfa", d => x"001bab"),
    (y => x"ede156", d => x"001ba4"),
    (y => x"edc5b7", d => x"001b9f"),
    (y => x"edaa20", d => x"001b97"),
    (y => x"ed8e8e", d => x"001b92"),
    (y => x"ed7303", d => x"001b8b"),
    (y => x"ed577f", d => x"001b84"),
    (y => x"ed3c01", d => x"001b7e"),
    (y => x"ed2089", d => x"001b78"),
    (y => x"ed0517", d => x"001b72"),
    (y => x"ece9ac", d => x"001b6b"),
    (y => x"ecce47", d => x"001b65"),
    (y => x"ecb2e9", d => x"001b5e"),
    (y => x"ec9791", d => x"001b58"),
    (y => x"ec7c3f", d => x"001b52"),
    (y => x"ec60f3", d => x"001b4c"),
    (y => x"ec45ae", d => x"001b45"),
    (y => x"ec2a6f", d => x"001b3f"),
    (y => x"ec0f37", d => x"001b38"),
    (y => x"ebf404", d => x"001b33"),
    (y => x"ebd8d8", d => x"001b2c"),
    (y => x"ebbdb2", d => x"001b26"),
    (y => x"eba293", d => x"001b1f"),
    (y => x"eb8779", d => x"001b1a"),
    (y => x"eb6c66", d => x"001b13"),
    (y => x"eb5159", d => x"001b0d"),
    (y => x"eb3653", d => x"001b06"),
    (y => x"eb1b52", d => x"001b01"),
    (y => x"eb0058", d => x"001afa"),
    (y => x"eae564", d => x"001af4"),
    (y => x"eaca76", d => x"001aee"),
    (y => x"eaaf8e", d => x"001ae8"),
    (y => x"ea94ac", d => x"001ae2"),
    (y => x"ea79d1", d => x"001adb"),
    (y => x"ea5efc", d => x"001ad5"),
    (y => x"ea442c", d => x"001ad0"),
    (y => x"ea2963", d => x"001ac9"),
    (y => x"ea0ea1", d => x"001ac2"),
    (y => x"e9f3e4", d => x"001abd"),
    (y => x"e9d92d", d => x"001ab7"),
    (y => x"e9be7c", d => x"001ab1"),
    (y => x"e9a3d2", d => x"001aaa"),
    (y => x"e9892e", d => x"001aa4"),
    (y => x"e96e8f", d => x"001a9f"),
    (y => x"e953f7", d => x"001a98"),
    (y => x"e93965", d => x"001a92"),
    (y => x"e91ed9", d => x"001a8c"),
    (y => x"e90452", d => x"001a87"),
    (y => x"e8e9d2", d => x"001a80"),
    (y => x"e8cf58", d => x"001a7a"),
    (y => x"e8b4e4", d => x"001a74"),
    (y => x"e89a76", d => x"001a6e"),
    (y => x"e8800e", d => x"001a68"),
    (y => x"e865ac", d => x"001a62"),
    (y => x"e84b50", d => x"001a5c"),
    (y => x"e830fa", d => x"001a56"),
    (y => x"e816aa", d => x"001a50"),
    (y => x"e7fc60", d => x"001a4a"),
    (y => x"e7e21b", d => x"001a45"),
    (y => x"e7c7dd", d => x"001a3e"),
    (y => x"e7ada5", d => x"001a38"),
    (y => x"e79373", d => x"001a32"),
    (y => x"e77946", d => x"001a2d"),
    (y => x"e75f1f", d => x"001a27"),
    (y => x"e744ff", d => x"001a20"),
    (y => x"e72ae4", d => x"001a1b"),
    (y => x"e710cf", d => x"001a15"),
    (y => x"e6f6c0", d => x"001a0f"),
    (y => x"e6dcb7", d => x"001a09"),
    (y => x"e6c2b4", d => x"001a03"),
    (y => x"e6a8b7", d => x"0019fd"),
    (y => x"e68ebf", d => x"0019f8"),
    (y => x"e674cd", d => x"0019f2"),
    (y => x"e65ae1", d => x"0019ec"),
    (y => x"e640fb", d => x"0019e6"),
    (y => x"e6271b", d => x"0019e0"),
    (y => x"e60d41", d => x"0019da"),
    (y => x"e5f36c", d => x"0019d5"),
    (y => x"e5d99e", d => x"0019ce"),
    (y => x"e5bfd5", d => x"0019c9"),
    (y => x"e5a611", d => x"0019c4"),
    (y => x"e58c54", d => x"0019bd"),
    (y => x"e5729c", d => x"0019b8"),
    (y => x"e558ea", d => x"0019b2"),
    (y => x"e53f3e", d => x"0019ac"),
    (y => x"e52598", d => x"0019a6"),
    (y => x"e50bf7", d => x"0019a1"),
    (y => x"e4f25c", d => x"00199b"),
    (y => x"e4d8c7", d => x"001995"),
    (y => x"e4bf37", d => x"001990"),
    (y => x"e4a5ae", d => x"001989"),
    (y => x"e48c2a", d => x"001984"),
    (y => x"e472ab", d => x"00197f"),
    (y => x"e45932", d => x"001979"),
    (y => x"e43fbf", d => x"001973"),
    (y => x"e42652", d => x"00196d"),
    (y => x"e40cea", d => x"001968"),
    (y => x"e3f388", d => x"001962"),
    (y => x"e3da2c", d => x"00195c"),
    (y => x"e3c0d5", d => x"001957"),
    (y => x"e3a784", d => x"001951"),
    (y => x"e38e39", d => x"00194b"),
    (y => x"e374f3", d => x"001946"),
    (y => x"e35bb2", d => x"001941"),
    (y => x"e34278", d => x"00193a"),
    (y => x"e32943", d => x"001935"),
    (y => x"e31013", d => x"001930"),
    (y => x"e2f6e9", d => x"00192a"),
    (y => x"e2ddc5", d => x"001924"),
    (y => x"e2c4a6", d => x"00191f"),
    (y => x"e2ab8d", d => x"001919"),
    (y => x"e29279", d => x"001914"),
    (y => x"e2796b", d => x"00190e"),
    (y => x"e26063", d => x"001908"),
    (y => x"e24760", d => x"001903"),
    (y => x"e22e62", d => x"0018fe"),
    (y => x"e2156a", d => x"0018f8"),
    (y => x"e1fc78", d => x"0018f2"),
    (y => x"e1e38b", d => x"0018ed"),
    (y => x"e1caa3", d => x"0018e8"),
    (y => x"e1b1c1", d => x"0018e2"),
    (y => x"e198e5", d => x"0018dc"),
    (y => x"e1800e", d => x"0018d7"),
    (y => x"e1673c", d => x"0018d2"),
    (y => x"e14e70", d => x"0018cc"),
    (y => x"e135a9", d => x"0018c7"),
    (y => x"e11ce8", d => x"0018c1"),
    (y => x"e1042c", d => x"0018bc"),
    (y => x"e0eb76", d => x"0018b6"),
    (y => x"e0d2c5", d => x"0018b1"),
    (y => x"e0ba1a", d => x"0018ab"),
    (y => x"e0a174", d => x"0018a6"),
    (y => x"e088d3", d => x"0018a1"),
    (y => x"e07038", d => x"00189b"),
    (y => x"e057a2", d => x"001896"),
    (y => x"e03f11", d => x"001891"),
    (y => x"e02686", d => x"00188b"),
    (y => x"e00e01", d => x"001885"),
    (y => x"dff580", d => x"001881"),
    (y => x"dfdd05", d => x"00187b"),
    (y => x"dfc48f", d => x"001876"),
    (y => x"dfac1f", d => x"001870"),
    (y => x"df93b4", d => x"00186b"),
    (y => x"df7b4e", d => x"001866"),
    (y => x"df62ee", d => x"001860"),
    (y => x"df4a93", d => x"00185b"),
    (y => x"df323d", d => x"001856"),
    (y => x"df19ed", d => x"001850"),
    (y => x"df01a2", d => x"00184b"),
    (y => x"dee95c", d => x"001846"),
    (y => x"ded11b", d => x"001841"),
    (y => x"deb8e0", d => x"00183b"),
    (y => x"dea0aa", d => x"001836"),
    (y => x"de8879", d => x"001831"),
    (y => x"de704e", d => x"00182b"),
    (y => x"de5828", d => x"001826"),
    (y => x"de4007", d => x"001821"),
    (y => x"de27eb", d => x"00181c"),
    (y => x"de0fd4", d => x"001817"),
    (y => x"ddf7c3", d => x"001811"),
    (y => x"dddfb7", d => x"00180c"),
    (y => x"ddc7b0", d => x"001807"),
    (y => x"ddafae", d => x"001802"),
    (y => x"dd97b2", d => x"0017fc"),
    (y => x"dd7fba", d => x"0017f8"),
    (y => x"dd67c8", d => x"0017f2"),
    (y => x"dd4fdb", d => x"0017ed"),
    (y => x"dd37f4", d => x"0017e7"),
    (y => x"dd2011", d => x"0017e3"),
    (y => x"dd0833", d => x"0017de"),
    (y => x"dcf05b", d => x"0017d8"),
    (y => x"dcd888", d => x"0017d3"),
    (y => x"dcc0ba", d => x"0017ce"),
    (y => x"dca8f1", d => x"0017c9"),
    (y => x"dc912d", d => x"0017c4"),
    (y => x"dc796f", d => x"0017be"),
    (y => x"dc61b5", d => x"0017ba"),
    (y => x"dc4a01", d => x"0017b4"),
    (y => x"dc3251", d => x"0017b0"),
    (y => x"dc1aa7", d => x"0017aa"),
    (y => x"dc0302", d => x"0017a5"),
    (y => x"dbeb62", d => x"0017a0"),
    (y => x"dbd3c7", d => x"00179b"),
    (y => x"dbbc31", d => x"001796"),
    (y => x"dba4a0", d => x"001791"),
    (y => x"db8d14", d => x"00178c"),
    (y => x"db758d", d => x"001787"),
    (y => x"db5e0b", d => x"001782"),
    (y => x"db468f", d => x"00177c"),
    (y => x"db2f17", d => x"001778"),
    (y => x"db17a4", d => x"001773"),
    (y => x"db0036", d => x"00176e"),
    (y => x"dae8ce", d => x"001768"),
    (y => x"dad16a", d => x"001764"),
    (y => x"daba0b", d => x"00175f"),
    (y => x"daa2b2", d => x"001759"),
    (y => x"da8b5d", d => x"001755"),
    (y => x"da740d", d => x"001750"),
    (y => x"da5cc3", d => x"00174a"),
    (y => x"da457d", d => x"001746"),
    (y => x"da2e3c", d => x"001741"),
    (y => x"da1700", d => x"00173c"),
    (y => x"d9ffc9", d => x"001737"),
    (y => x"d9e897", d => x"001732"),
    (y => x"d9d16a", d => x"00172d"),
    (y => x"d9ba42", d => x"001728"),
    (y => x"d9a31f", d => x"001723"),
    (y => x"d98c01", d => x"00171e"),
    (y => x"d974e7", d => x"00171a"),
    (y => x"d95dd3", d => x"001714"),
    (y => x"d946c3", d => x"001710"),
    (y => x"d92fb8", d => x"00170b"),
    (y => x"d918b3", d => x"001705"),
    (y => x"d901b2", d => x"001701"),
    (y => x"d8eab6", d => x"0016fc"),
    (y => x"d8d3be", d => x"0016f8"),
    (y => x"d8bccc", d => x"0016f2"),
    (y => x"d8a5df", d => x"0016ed"),
    (y => x"d88ef6", d => x"0016e9"),
    (y => x"d87812", d => x"0016e4"),
    (y => x"d86133", d => x"0016df"),
    (y => x"d84a59", d => x"0016da"),
    (y => x"d83384", d => x"0016d5"),
    (y => x"d81cb4", d => x"0016d0"),
    (y => x"d805e8", d => x"0016cc"),
    (y => x"d7ef21", d => x"0016c7"),
    (y => x"d7d85f", d => x"0016c2"),
    (y => x"d7c1a2", d => x"0016bd"),
    (y => x"d7aae9", d => x"0016b9"),
    (y => x"d79436", d => x"0016b3"),
    (y => x"d77d87", d => x"0016af"),
    (y => x"d766dd", d => x"0016aa"),
    (y => x"d75037", d => x"0016a6"),
    (y => x"d73997", d => x"0016a0"),
    (y => x"d722fb", d => x"00169c"),
    (y => x"d70c64", d => x"001697"),
    (y => x"d6f5d1", d => x"001693"),
    (y => x"d6df44", d => x"00168d"),
    (y => x"d6c8bb", d => x"001689"),
    (y => x"d6b237", d => x"001684"),
    (y => x"d69bb7", d => x"001680"),
    (y => x"d6853c", d => x"00167b"),
    (y => x"d66ec6", d => x"001676"),
    (y => x"d65855", d => x"001671"),
    (y => x"d641e8", d => x"00166d"),
    (y => x"d62b81", d => x"001667"),
    (y => x"d6151d", d => x"001664"),
    (y => x"d5febf", d => x"00165e"),
    (y => x"d5e865", d => x"00165a"),
    (y => x"d5d210", d => x"001655"),
    (y => x"d5bbbf", d => x"001651"),
    (y => x"d5a573", d => x"00164c"),
    (y => x"d58f2c", d => x"001647"),
    (y => x"d578e9", d => x"001643"),
    (y => x"d562ab", d => x"00163e"),
    (y => x"d54c72", d => x"001639"),
    (y => x"d5363d", d => x"001635"),
    (y => x"d5200d", d => x"001630"),
    (y => x"d509e2", d => x"00162b"),
    (y => x"d4f3bb", d => x"001627"),
    (y => x"d4dd98", d => x"001623"),
    (y => x"d4c77b", d => x"00161d"),
    (y => x"d4b162", d => x"001619"),
    (y => x"d49b4d", d => x"001615"),
    (y => x"d4853d", d => x"001610"),
    (y => x"d46f32", d => x"00160b"),
    (y => x"d4592b", d => x"001607"),
    (y => x"d44329", d => x"001602"),
    (y => x"d42d2b", d => x"0015fe"),
    (y => x"d41732", d => x"0015f9"),
    (y => x"d4013e", d => x"0015f4"),
    (y => x"d3eb4e", d => x"0015f0"),
    (y => x"d3d562", d => x"0015ec"),
    (y => x"d3bf7b", d => x"0015e7"),
    (y => x"d3a999", d => x"0015e2"),
    (y => x"d393bb", d => x"0015de"),
    (y => x"d37de2", d => x"0015d9"),
    (y => x"d3680d", d => x"0015d5"),
    (y => x"d3523d", d => x"0015d0"),
    (y => x"d33c71", d => x"0015cc"),
    (y => x"d326a9", d => x"0015c8"),
    (y => x"d310e7", d => x"0015c2"),
    (y => x"d2fb28", d => x"0015bf"),
    (y => x"d2e56e", d => x"0015ba"),
    (y => x"d2cfb9", d => x"0015b5"),
    (y => x"d2ba08", d => x"0015b1"),
    (y => x"d2a45b", d => x"0015ad"),
    (y => x"d28eb3", d => x"0015a8"),
    (y => x"d27910", d => x"0015a3"),
    (y => x"d26371", d => x"00159f"),
    (y => x"d24dd6", d => x"00159b"),
    (y => x"d23840", d => x"001596"),
    (y => x"d222ae", d => x"001592"),
    (y => x"d20d21", d => x"00158d"),
    (y => x"d1f798", d => x"001589"),
    (y => x"d1e213", d => x"001585"),
    (y => x"d1cc93", d => x"001580"),
    (y => x"d1b717", d => x"00157c"),
    (y => x"d1a1a0", d => x"001577"),
    (y => x"d18c2d", d => x"001573"),
    (y => x"d176be", d => x"00156f"),
    (y => x"d16154", d => x"00156a"),
    (y => x"d14bee", d => x"001566"),
    (y => x"d1368d", d => x"001561"),
    (y => x"d12130", d => x"00155d"),
    (y => x"d10bd7", d => x"001559"),
    (y => x"d0f683", d => x"001554"),
    (y => x"d0e133", d => x"001550"),
    (y => x"d0cbe7", d => x"00154c"),
    (y => x"d0b6a0", d => x"001547"),
    (y => x"d0a15d", d => x"001543"),
    (y => x"d08c1e", d => x"00153f"),
    (y => x"d076e4", d => x"00153a"),
    (y => x"d061ae", d => x"001536"),
    (y => x"d04c7c", d => x"001532"),
    (y => x"d0374e", d => x"00152e"),
    (y => x"d02225", d => x"001529"),
    (y => x"d00d01", d => x"001524"),
    (y => x"cff7e0", d => x"001521"),
    (y => x"cfe2c4", d => x"00151c"),
    (y => x"cfcdac", d => x"001518"),
    (y => x"cfb898", d => x"001514"),
    (y => x"cfa389", d => x"00150f"),
    (y => x"cf8e7e", d => x"00150b"),
    (y => x"cf7977", d => x"001507"),
    (y => x"cf6474", d => x"001503"),
    (y => x"cf4f76", d => x"0014fe"),
    (y => x"cf3a7c", d => x"0014fa"),
    (y => x"cf2586", d => x"0014f6"),
    (y => x"cf1095", d => x"0014f1"),
    (y => x"cefba7", d => x"0014ee"),
    (y => x"cee6be", d => x"0014e9"),
    (y => x"ced1d9", d => x"0014e5"),
    (y => x"cebcf8", d => x"0014e1"),
    (y => x"cea81c", d => x"0014dc"),
    (y => x"ce9344", d => x"0014d8"),
    (y => x"ce7e70", d => x"0014d4"),
    (y => x"ce69a0", d => x"0014d0"),
    (y => x"ce54d4", d => x"0014cc"),
    (y => x"ce400d", d => x"0014c7"),
    (y => x"ce2b49", d => x"0014c4"),
    (y => x"ce168a", d => x"0014bf"),
    (y => x"ce01cf", d => x"0014bb"),
    (y => x"cded18", d => x"0014b7"),
    (y => x"cdd866", d => x"0014b2"),
    (y => x"cdc3b7", d => x"0014af"),
    (y => x"cdaf0d", d => x"0014aa"),
    (y => x"cd9a67", d => x"0014a6"),
    (y => x"cd85c5", d => x"0014a2"),
    (y => x"cd7127", d => x"00149e"),
    (y => x"cd5c8d", d => x"00149a"),
    (y => x"cd47f8", d => x"001495"),
    (y => x"cd3366", d => x"001492"),
    (y => x"cd1ed9", d => x"00148d"),
    (y => x"cd0a50", d => x"001489"),
    (y => x"ccf5cb", d => x"001485"),
    (y => x"cce149", d => x"001482"),
    (y => x"cccccd", d => x"00147c"),
    (y => x"ccb854", d => x"001479"),
    (y => x"cca3df", d => x"001475"),
    (y => x"cc8f6e", d => x"001471"),
    (y => x"cc7b02", d => x"00146c"),
    (y => x"cc6699", d => x"001469"),
    (y => x"cc5235", d => x"001464"),
    (y => x"cc3dd4", d => x"001461"),
    (y => x"cc2978", d => x"00145c"),
    (y => x"cc1520", d => x"001458"),
    (y => x"cc00cc", d => x"001454"),
    (y => x"cbec7c", d => x"001450"),
    (y => x"cbd830", d => x"00144c"),
    (y => x"cbc3e7", d => x"001449"),
    (y => x"cbafa3", d => x"001444"),
    (y => x"cb9b63", d => x"001440"),
    (y => x"cb8728", d => x"00143b"),
    (y => x"cb72f0", d => x"001438"),
    (y => x"cb5ebc", d => x"001434"),
    (y => x"cb4a8c", d => x"001430"),
    (y => x"cb3660", d => x"00142c"),
    (y => x"cb2238", d => x"001428"),
    (y => x"cb0e14", d => x"001424"),
    (y => x"caf9f4", d => x"001420"),
    (y => x"cae5d8", d => x"00141c"),
    (y => x"cad1c0", d => x"001418"),
    (y => x"cabdac", d => x"001414"),
    (y => x"caa99c", d => x"001410"),
    (y => x"ca9590", d => x"00140c"),
    (y => x"ca8188", d => x"001408"),
    (y => x"ca6d84", d => x"001404"),
    (y => x"ca5984", d => x"001400"),
    (y => x"ca4588", d => x"0013fc"),
    (y => x"ca318f", d => x"0013f9"),
    (y => x"ca1d9b", d => x"0013f4"),
    (y => x"ca09ab", d => x"0013f0"),
    (y => x"c9f5be", d => x"0013ed"),
    (y => x"c9e1d6", d => x"0013e8"),
    (y => x"c9cdf1", d => x"0013e5"),
    (y => x"c9ba11", d => x"0013e0"),
    (y => x"c9a634", d => x"0013dd"),
    (y => x"c9925b", d => x"0013d9"),
    (y => x"c97e86", d => x"0013d5"),
    (y => x"c96ab5", d => x"0013d1"),
    (y => x"c956e8", d => x"0013cd"),
    (y => x"c9431f", d => x"0013c9"),
    (y => x"c92f59", d => x"0013c6"),
    (y => x"c91b98", d => x"0013c1"),
    (y => x"c907da", d => x"0013be"),
    (y => x"c8f420", d => x"0013ba"),
    (y => x"c8e06a", d => x"0013b6"),
    (y => x"c8ccb8", d => x"0013b2"),
    (y => x"c8b90a", d => x"0013ae"),
    (y => x"c8a560", d => x"0013aa"),
    (y => x"c891ba", d => x"0013a6"),
    (y => x"c87e17", d => x"0013a3"),
    (y => x"c86a78", d => x"00139f"),
    (y => x"c856dd", d => x"00139b"),
    (y => x"c84346", d => x"001397"),
    (y => x"c82fb3", d => x"001393"),
    (y => x"c81c24", d => x"00138f"),
    (y => x"c80898", d => x"00138c"),
    (y => x"c7f510", d => x"001388"),
    (y => x"c7e18c", d => x"001384"),
    (y => x"c7ce0c", d => x"001380"),
    (y => x"c7ba90", d => x"00137c"),
    (y => x"c7a717", d => x"001379"),
    (y => x"c793a3", d => x"001374"),
    (y => x"c78032", d => x"001371"),
    (y => x"c76cc4", d => x"00136e"),
    (y => x"c7595b", d => x"001369"),
    (y => x"c745f5", d => x"001366"),
    (y => x"c73294", d => x"001361"),
    (y => x"c71f36", d => x"00135e"),
    (y => x"c70bdb", d => x"00135b"),
    (y => x"c6f885", d => x"001356"),
    (y => x"c6e532", d => x"001353"),
    (y => x"c6d1e3", d => x"00134f"),
    (y => x"c6be98", d => x"00134b"),
    (y => x"c6ab50", d => x"001348"),
    (y => x"c6980c", d => x"001344"),
    (y => x"c684cc", d => x"001340"),
    (y => x"c67190", d => x"00133c"),
    (y => x"c65e57", d => x"001339"),
    (y => x"c64b22", d => x"001335"),
    (y => x"c637f1", d => x"001331"),
    (y => x"c624c4", d => x"00132d"),
    (y => x"c6119a", d => x"00132a"),
    (y => x"c5fe74", d => x"001326"),
    (y => x"c5eb51", d => x"001323"),
    (y => x"c5d833", d => x"00131e"),
    (y => x"c5c518", d => x"00131b"),
    (y => x"c5b201", d => x"001317"),
    (y => x"c59eed", d => x"001314"),
    (y => x"c58bdd", d => x"001310"),
    (y => x"c578d1", d => x"00130c"),
    (y => x"c565c8", d => x"001309"),
    (y => x"c552c3", d => x"001305"),
    (y => x"c53fc2", d => x"001301"),
    (y => x"c52cc5", d => x"0012fd"),
    (y => x"c519cb", d => x"0012fa"),
    (y => x"c506d4", d => x"0012f7"),
    (y => x"c4f3e2", d => x"0012f2"),
    (y => x"c4e0f3", d => x"0012ef"),
    (y => x"c4ce07", d => x"0012ec"),
    (y => x"c4bb20", d => x"0012e7"),
    (y => x"c4a83c", d => x"0012e4"),
    (y => x"c4955b", d => x"0012e1"),
    (y => x"c4827e", d => x"0012dd"),
    (y => x"c46fa5", d => x"0012d9"),
    (y => x"c45cd0", d => x"0012d5"),
    (y => x"c449fe", d => x"0012d2"),
    (y => x"c4372f", d => x"0012cf"),
    (y => x"c42465", d => x"0012ca"),
    (y => x"c4119d", d => x"0012c8"),
    (y => x"c3feda", d => x"0012c3"),
    (y => x"c3ec1a", d => x"0012c0"),
    (y => x"c3d95d", d => x"0012bd"),
    (y => x"c3c6a5", d => x"0012b8"),
    (y => x"c3b3ef", d => x"0012b6"),
    (y => x"c3a13e", d => x"0012b1"),
    (y => x"c38e90", d => x"0012ae"),
    (y => x"c37be5", d => x"0012ab"),
    (y => x"c3693e", d => x"0012a7"),
    (y => x"c3569b", d => x"0012a3"),
    (y => x"c343fb", d => x"0012a0"),
    (y => x"c3315f", d => x"00129c"),
    (y => x"c31ec6", d => x"001299"),
    (y => x"c30c31", d => x"001295"),
    (y => x"c2f99f", d => x"001292"),
    (y => x"c2e711", d => x"00128e"),
    (y => x"c2d486", d => x"00128b"),
    (y => x"c2c1ff", d => x"001287"),
    (y => x"c2af7b", d => x"001284"),
    (y => x"c29cfb", d => x"001280"),
    (y => x"c28a7f", d => x"00127c"),
    (y => x"c27806", d => x"001279"),
    (y => x"c26590", d => x"001276"),
    (y => x"c2531e", d => x"001272"),
    (y => x"c240b0", d => x"00126e"),
    (y => x"c22e45", d => x"00126b"),
    (y => x"c21bdd", d => x"001268"),
    (y => x"c20979", d => x"001264"),
    (y => x"c1f719", d => x"001260"),
    (y => x"c1e4bc", d => x"00125d"),
    (y => x"c1d262", d => x"00125a"),
    (y => x"c1c00c", d => x"001256"),
    (y => x"c1adb9", d => x"001253"),
    (y => x"c19b6a", d => x"00124f"),
    (y => x"c1891e", d => x"00124c"),
    (y => x"c176d6", d => x"001248"),
    (y => x"c16491", d => x"001245"),
    (y => x"c15250", d => x"001241"),
    (y => x"c14012", d => x"00123e"),
    (y => x"c12dd7", d => x"00123b"),
    (y => x"c11ba0", d => x"001237"),
    (y => x"c1096d", d => x"001233"),
    (y => x"c0f73d", d => x"001230"),
    (y => x"c0e510", d => x"00122d"),
    (y => x"c0d2e6", d => x"00122a"),
    (y => x"c0c0c1", d => x"001225"),
    (y => x"c0ae9e", d => x"001223"),
    (y => x"c09c7f", d => x"00121f"),
    (y => x"c08a63", d => x"00121c"),
    (y => x"c0784b", d => x"001218"),
    (y => x"c06636", d => x"001215"),
    (y => x"c05425", d => x"001211"),
    (y => x"c04217", d => x"00120e"),
    (y => x"c0300c", d => x"00120b"),
    (y => x"c01e04", d => x"001208"),
    (y => x"c00c01", d => x"001203"),
    (y => x"bffa00", d => x"001201"),
    (y => x"bfe803", d => x"0011fd"),
    (y => x"bfd609", d => x"0011fa"),
    (y => x"bfc413", d => x"0011f6"),
    (y => x"bfb21f", d => x"0011f4"),
    (y => x"bfa030", d => x"0011ef"),
    (y => x"bf8e43", d => x"0011ed"),
    (y => x"bf7c5a", d => x"0011e9"),
    (y => x"bf6a75", d => x"0011e5"),
    (y => x"bf5892", d => x"0011e3"),
    (y => x"bf46b3", d => x"0011df"),
    (y => x"bf34d8", d => x"0011db"),
    (y => x"bf22ff", d => x"0011d9"),
    (y => x"bf112a", d => x"0011d5"),
    (y => x"beff59", d => x"0011d1"),
    (y => x"beed8a", d => x"0011cf"),
    (y => x"bedbbf", d => x"0011cb"),
    (y => x"bec9f8", d => x"0011c7"),
    (y => x"beb833", d => x"0011c5"),
    (y => x"bea672", d => x"0011c1"),
    (y => x"be94b4", d => x"0011be"),
    (y => x"be82fa", d => x"0011ba"),
    (y => x"be7143", d => x"0011b7"),
    (y => x"be5f8f", d => x"0011b4"),
    (y => x"be4dde", d => x"0011b1"),
    (y => x"be3c31", d => x"0011ad"),
    (y => x"be2a87", d => x"0011aa"),
    (y => x"be18e0", d => x"0011a7"),
    (y => x"be073d", d => x"0011a3"),
    (y => x"bdf59c", d => x"0011a1"),
    (y => x"bde3ff", d => x"00119d"),
    (y => x"bdd266", d => x"001199"),
    (y => x"bdc0cf", d => x"001197"),
    (y => x"bdaf3c", d => x"001193"),
    (y => x"bd9dac", d => x"001190"),
    (y => x"bd8c20", d => x"00118c"),
    (y => x"bd7a96", d => x"00118a"),
    (y => x"bd6910", d => x"001186"),
    (y => x"bd578d", d => x"001183"),
    (y => x"bd460d", d => x"001180"),
    (y => x"bd3491", d => x"00117c"),
    (y => x"bd2318", d => x"001179"),
    (y => x"bd11a2", d => x"001176"),
    (y => x"bd002f", d => x"001173"),
    (y => x"bceebf", d => x"001170"),
    (y => x"bcdd53", d => x"00116c"),
    (y => x"bccbea", d => x"001169"),
    (y => x"bcba84", d => x"001166"),
    (y => x"bca921", d => x"001163"),
    (y => x"bc97c2", d => x"00115f"),
    (y => x"bc8666", d => x"00115c"),
    (y => x"bc750c", d => x"00115a"),
    (y => x"bc63b7", d => x"001155"),
    (y => x"bc5264", d => x"001153"),
    (y => x"bc4114", d => x"001150"),
    (y => x"bc2fc8", d => x"00114c"),
    (y => x"bc1e7f", d => x"001149"),
    (y => x"bc0d39", d => x"001146"),
    (y => x"bbfbf6", d => x"001143"),
    (y => x"bbeab6", d => x"001140"),
    (y => x"bbd97a", d => x"00113c"),
    (y => x"bbc840", d => x"00113a"),
    (y => x"bbb70a", d => x"001136"),
    (y => x"bba5d7", d => x"001133"),
    (y => x"bb94a7", d => x"001130"),
    (y => x"bb837a", d => x"00112d"),
    (y => x"bb7251", d => x"001129"),
    (y => x"bb612a", d => x"001127"),
    (y => x"bb5007", d => x"001123"),
    (y => x"bb3ee7", d => x"001120"),
    (y => x"bb2dca", d => x"00111d"),
    (y => x"bb1cb0", d => x"00111a"),
    (y => x"bb0b99", d => x"001117"),
    (y => x"bafa85", d => x"001114"),
    (y => x"bae975", d => x"001110"),
    (y => x"bad867", d => x"00110e"),
    (y => x"bac75d", d => x"00110a"),
    (y => x"bab656", d => x"001107"),
    (y => x"baa552", d => x"001104"),
    (y => x"ba9451", d => x"001101"),
    (y => x"ba8353", d => x"0010fe"),
    (y => x"ba7258", d => x"0010fb"),
    (y => x"ba6160", d => x"0010f8"),
    (y => x"ba506c", d => x"0010f4"),
    (y => x"ba3f7a", d => x"0010f2"),
    (y => x"ba2e8b", d => x"0010ef"),
    (y => x"ba1da0", d => x"0010eb"),
    (y => x"ba0cb8", d => x"0010e8"),
    (y => x"b9fbd2", d => x"0010e6"),
    (y => x"b9eaf0", d => x"0010e2"),
    (y => x"b9da11", d => x"0010df"),
    (y => x"b9c935", d => x"0010dc"),
    (y => x"b9b85c", d => x"0010d9"),
    (y => x"b9a786", d => x"0010d6"),
    (y => x"b996b3", d => x"0010d3"),
    (y => x"b985e3", d => x"0010d0"),
    (y => x"b97516", d => x"0010cd"),
    (y => x"b9644d", d => x"0010c9"),
    (y => x"b95386", d => x"0010c7"),
    (y => x"b942c2", d => x"0010c4"),
    (y => x"b93201", d => x"0010c1"),
    (y => x"b92144", d => x"0010bd"),
    (y => x"b91089", d => x"0010bb"),
    (y => x"b8ffd2", d => x"0010b7"),
    (y => x"b8ef1d", d => x"0010b5"),
    (y => x"b8de6b", d => x"0010b2"),
    (y => x"b8cdbd", d => x"0010ae"),
    (y => x"b8bd11", d => x"0010ac"),
    (y => x"b8ac69", d => x"0010a8"),
    (y => x"b89bc3", d => x"0010a6"),
    (y => x"b88b21", d => x"0010a2"),
    (y => x"b87a81", d => x"0010a0"),
    (y => x"b869e5", d => x"00109c"),
    (y => x"b8594b", d => x"00109a"),
    (y => x"b848b4", d => x"001097"),
    (y => x"b83821", d => x"001093"),
    (y => x"b82790", d => x"001091"),
    (y => x"b81703", d => x"00108d"),
    (y => x"b80678", d => x"00108b"),
    (y => x"b7f5f0", d => x"001088"),
    (y => x"b7e56c", d => x"001084"),
    (y => x"b7d4ea", d => x"001082"),
    (y => x"b7c46b", d => x"00107f"),
    (y => x"b7b3ef", d => x"00107c"),
    (y => x"b7a376", d => x"001079"),
    (y => x"b79301", d => x"001075"),
    (y => x"b7828e", d => x"001073"),
    (y => x"b7721e", d => x"001070"),
    (y => x"b761b0", d => x"00106e"),
    (y => x"b75146", d => x"00106a"),
    (y => x"b740df", d => x"001067"),
    (y => x"b7307b", d => x"001064"),
    (y => x"b7201a", d => x"001061"),
    (y => x"b70fbb", d => x"00105f"),
    (y => x"b6ff60", d => x"00105b"),
    (y => x"b6ef07", d => x"001059"),
    (y => x"b6deb2", d => x"001055"),
    (y => x"b6ce5f", d => x"001053"),
    (y => x"b6be0f", d => x"001050"),
    (y => x"b6adc2", d => x"00104d"),
    (y => x"b69d78", d => x"00104a"),
    (y => x"b68d31", d => x"001047"),
    (y => x"b67ced", d => x"001044"),
    (y => x"b66cac", d => x"001041"),
    (y => x"b65c6d", d => x"00103f"),
    (y => x"b64c32", d => x"00103b"),
    (y => x"b63bf9", d => x"001039"),
    (y => x"b62bc3", d => x"001036"),
    (y => x"b61b90", d => x"001033"),
    (y => x"b60b61", d => x"00102f"),
    (y => x"b5fb33", d => x"00102e"),
    (y => x"b5eb09", d => x"00102a"),
    (y => x"b5dae2", d => x"001027"),
    (y => x"b5cabd", d => x"001025"),
    (y => x"b5ba9c", d => x"001021"),
    (y => x"b5aa7d", d => x"00101f"),
    (y => x"b59a61", d => x"00101c"),
    (y => x"b58a48", d => x"001019"),
    (y => x"b57a32", d => x"001016"),
    (y => x"b56a1f", d => x"001013"),
    (y => x"b55a0e", d => x"001011"),
    (y => x"b54a01", d => x"00100d"),
    (y => x"b539f6", d => x"00100b"),
    (y => x"b529ee", d => x"001008"),
    (y => x"b519e9", d => x"001005"),
    (y => x"b509e6", d => x"001003"),
    (y => x"b4f9e7", d => x"000fff"),
    (y => x"b4e9ea", d => x"000ffd"),
    (y => x"b4d9f0", d => x"000ffa"),
    (y => x"b4c9f9", d => x"000ff7"),
    (y => x"b4ba05", d => x"000ff4"),
    (y => x"b4aa14", d => x"000ff1"),
    (y => x"b49a25", d => x"000fef"),
    (y => x"b48a3a", d => x"000feb"),
    (y => x"b47a51", d => x"000fe9"),
    (y => x"b46a6b", d => x"000fe6"),
    (y => x"b45a87", d => x"000fe4"),
    (y => x"b44aa7", d => x"000fe0"),
    (y => x"b43ac9", d => x"000fde"),
    (y => x"b42aee", d => x"000fdb"),
    (y => x"b41b16", d => x"000fd8"),
    (y => x"b40b41", d => x"000fd5"),
    (y => x"b3fb6e", d => x"000fd3"),
    (y => x"b3eb9e", d => x"000fd0"),
    (y => x"b3dbd1", d => x"000fcd"),
    (y => x"b3cc07", d => x"000fca"),
    (y => x"b3bc3f", d => x"000fc8"),
    (y => x"b3ac7b", d => x"000fc4"),
    (y => x"b39cb9", d => x"000fc2"),
    (y => x"b38cfa", d => x"000fbf"),
    (y => x"b37d3d", d => x"000fbd"),
    (y => x"b36d83", d => x"000fba"),
    (y => x"b35dcd", d => x"000fb6"),
    (y => x"b34e18", d => x"000fb5"),
    (y => x"b33e67", d => x"000fb1"),
    (y => x"b32eb8", d => x"000faf"),
    (y => x"b31f0c", d => x"000fac"),
    (y => x"b30f63", d => x"000fa9"),
    (y => x"b2ffbd", d => x"000fa6"),
    (y => x"b2f019", d => x"000fa4"),
    (y => x"b2e078", d => x"000fa1"),
    (y => x"b2d0da", d => x"000f9e"),
    (y => x"b2c13e", d => x"000f9c"),
    (y => x"b2b1a5", d => x"000f99"),
    (y => x"b2a20f", d => x"000f96"),
    (y => x"b2927c", d => x"000f93"),
    (y => x"b282eb", d => x"000f91"),
    (y => x"b2735d", d => x"000f8e"),
    (y => x"b263d2", d => x"000f8b"),
    (y => x"b2544a", d => x"000f88"),
    (y => x"b244c4", d => x"000f86"),
    (y => x"b23541", d => x"000f83"),
    (y => x"b225c0", d => x"000f81"),
    (y => x"b21643", d => x"000f7d"),
    (y => x"b206c8", d => x"000f7b"),
    (y => x"b1f74f", d => x"000f79"),
    (y => x"b1e7da", d => x"000f75"),
    (y => x"b1d867", d => x"000f73"),
    (y => x"b1c8f6", d => x"000f71"),
    (y => x"b1b989", d => x"000f6d"),
    (y => x"b1aa1e", d => x"000f6b"),
    (y => x"b19ab6", d => x"000f68"),
    (y => x"b18b50", d => x"000f66"),
    (y => x"b17bed", d => x"000f63"),
    (y => x"b16c8d", d => x"000f60"),
    (y => x"b15d2f", d => x"000f5e"),
    (y => x"b14dd4", d => x"000f5b"),
    (y => x"b13e7c", d => x"000f58"),
    (y => x"b12f27", d => x"000f55"),
    (y => x"b11fd4", d => x"000f53"),
    (y => x"b11083", d => x"000f51"),
    (y => x"b10136", d => x"000f4d"),
    (y => x"b0f1eb", d => x"000f4b"),
    (y => x"b0e2a2", d => x"000f49"),
    (y => x"b0d35c", d => x"000f46"),
    (y => x"b0c419", d => x"000f43"),
    (y => x"b0b4d9", d => x"000f40"),
    (y => x"b0a59b", d => x"000f3e"),
    (y => x"b09660", d => x"000f3b"),
    (y => x"b08727", d => x"000f39"),
    (y => x"b077f1", d => x"000f36"),
    (y => x"b068be", d => x"000f33"),
    (y => x"b0598d", d => x"000f31"),
    (y => x"b04a5f", d => x"000f2e"),
    (y => x"b03b34", d => x"000f2b"),
    (y => x"b02c0b", d => x"000f29"),
    (y => x"b01ce5", d => x"000f26"),
    (y => x"b00dc1", d => x"000f24"),
    (y => x"affea0", d => x"000f21"),
    (y => x"afef81", d => x"000f1f"),
    (y => x"afe066", d => x"000f1b"),
    (y => x"afd14c", d => x"000f1a"),
    (y => x"afc236", d => x"000f16"),
    (y => x"afb321", d => x"000f15"),
    (y => x"afa410", d => x"000f11"),
    (y => x"af9501", d => x"000f0f"),
    (y => x"af85f5", d => x"000f0c"),
    (y => x"af76eb", d => x"000f0a"),
    (y => x"af67e4", d => x"000f07"),
    (y => x"af58df", d => x"000f05"),
    (y => x"af49dd", d => x"000f02"),
    (y => x"af3ade", d => x"000eff"),
    (y => x"af2be1", d => x"000efd"),
    (y => x"af1ce6", d => x"000efb"),
    (y => x"af0def", d => x"000ef7"),
    (y => x"aefef9", d => x"000ef6"),
    (y => x"aef007", d => x"000ef2"),
    (y => x"aee117", d => x"000ef0"),
    (y => x"aed229", d => x"000eee"),
    (y => x"aec33e", d => x"000eeb"),
    (y => x"aeb455", d => x"000ee9"),
    (y => x"aea570", d => x"000ee5"),
    (y => x"ae968c", d => x"000ee4"),
    (y => x"ae87ab", d => x"000ee1"),
    (y => x"ae78cd", d => x"000ede"),
    (y => x"ae69f1", d => x"000edc"),
    (y => x"ae5b18", d => x"000ed9"),
    (y => x"ae4c41", d => x"000ed7"),
    (y => x"ae3d6d", d => x"000ed4"),
    (y => x"ae2e9b", d => x"000ed2"),
    (y => x"ae1fcc", d => x"000ecf"),
    (y => x"ae1100", d => x"000ecc"),
    (y => x"ae0235", d => x"000ecb"),
    (y => x"adf36e", d => x"000ec7"),
    (y => x"ade4a9", d => x"000ec5"),
    (y => x"add5e6", d => x"000ec3"),
    (y => x"adc726", d => x"000ec0"),
    (y => x"adb868", d => x"000ebe"),
    (y => x"ada9ad", d => x"000ebb"),
    (y => x"ad9af5", d => x"000eb8"),
    (y => x"ad8c3f", d => x"000eb6"),
    (y => x"ad7d8b", d => x"000eb4"),
    (y => x"ad6eda", d => x"000eb1"),
    (y => x"ad602b", d => x"000eaf"),
    (y => x"ad517f", d => x"000eac"),
    (y => x"ad42d5", d => x"000eaa"),
    (y => x"ad342e", d => x"000ea7"),
    (y => x"ad2589", d => x"000ea5"),
    (y => x"ad16e7", d => x"000ea2"),
    (y => x"ad0847", d => x"000ea0"),
    (y => x"acf9aa", d => x"000e9d"),
    (y => x"aceb0f", d => x"000e9b"),
    (y => x"acdc77", d => x"000e98"),
    (y => x"accde1", d => x"000e96"),
    (y => x"acbf4e", d => x"000e93"),
    (y => x"acb0bd", d => x"000e91"),
    (y => x"aca22e", d => x"000e8f"),
    (y => x"ac93a2", d => x"000e8c"),
    (y => x"ac8519", d => x"000e89"),
    (y => x"ac7691", d => x"000e88"),
    (y => x"ac680d", d => x"000e84"),
    (y => x"ac598a", d => x"000e83"),
    (y => x"ac4b0b", d => x"000e7f"),
    (y => x"ac3c8d", d => x"000e7e"),
    (y => x"ac2e12", d => x"000e7b"),
    (y => x"ac1f9a", d => x"000e78"),
    (y => x"ac1124", d => x"000e76"),
    (y => x"ac02b0", d => x"000e74"),
    (y => x"abf43f", d => x"000e71"),
    (y => x"abe5d0", d => x"000e6f"),
    (y => x"abd763", d => x"000e6d"),
    (y => x"abc8f9", d => x"000e6a"),
    (y => x"abba92", d => x"000e67"),
    (y => x"abac2d", d => x"000e65"),
    (y => x"ab9dca", d => x"000e63"),
    (y => x"ab8f6a", d => x"000e60"),
    (y => x"ab810c", d => x"000e5e"),
    (y => x"ab72b0", d => x"000e5c"),
    (y => x"ab6457", d => x"000e59"),
    (y => x"ab5601", d => x"000e56"),
    (y => x"ab47ac", d => x"000e55"),
    (y => x"ab395a", d => x"000e52"),
    (y => x"ab2b0b", d => x"000e4f"),
    (y => x"ab1cbe", d => x"000e4d"),
    (y => x"ab0e73", d => x"000e4b"),
    (y => x"ab002b", d => x"000e48"),
    (y => x"aaf1e5", d => x"000e46"),
    (y => x"aae3a1", d => x"000e44"),
    (y => x"aad560", d => x"000e41"),
    (y => x"aac721", d => x"000e3f"),
    (y => x"aab8e5", d => x"000e3c"),
    (y => x"aaaaab", d => x"000e3a"),
    (y => x"aa9c73", d => x"000e38"),
    (y => x"aa8e3d", d => x"000e36"),
    (y => x"aa800b", d => x"000e32"),
    (y => x"aa71da", d => x"000e31"),
    (y => x"aa63ac", d => x"000e2e"),
    (y => x"aa5580", d => x"000e2c"),
    (y => x"aa4756", d => x"000e2a"),
    (y => x"aa392f", d => x"000e27"),
    (y => x"aa2b0a", d => x"000e25"),
    (y => x"aa1ce8", d => x"000e22"),
    (y => x"aa0ec8", d => x"000e20"),
    (y => x"aa00aa", d => x"000e1e"),
    (y => x"a9f28e", d => x"000e1c"),
    (y => x"a9e475", d => x"000e19"),
    (y => x"a9d65f", d => x"000e16"),
    (y => x"a9c84a", d => x"000e15"),
    (y => x"a9ba38", d => x"000e12"),
    (y => x"a9ac28", d => x"000e10"),
    (y => x"a99e1b", d => x"000e0d"),
    (y => x"a99010", d => x"000e0b"),
    (y => x"a98207", d => x"000e09"),
    (y => x"a97401", d => x"000e06"),
    (y => x"a965fc", d => x"000e05"),
    (y => x"a957fb", d => x"000e01"),
    (y => x"a949fb", d => x"000e00"),
    (y => x"a93bfe", d => x"000dfd"),
    (y => x"a92e03", d => x"000dfb"),
    (y => x"a9200a", d => x"000df9"),
    (y => x"a91214", d => x"000df6"),
    (y => x"a90420", d => x"000df4"),
    (y => x"a8f62f", d => x"000df1"),
    (y => x"a8e83f", d => x"000df0"),
    (y => x"a8da52", d => x"000ded"),
    (y => x"a8cc67", d => x"000deb"),
    (y => x"a8be7f", d => x"000de8"),
    (y => x"a8b099", d => x"000de6"),
    (y => x"a8a2b5", d => x"000de4"),
    (y => x"a894d3", d => x"000de2"),
    (y => x"a886f4", d => x"000ddf"),
    (y => x"a87917", d => x"000ddd"),
    (y => x"a86b3c", d => x"000ddb"),
    (y => x"a85d64", d => x"000dd8"),
    (y => x"a84f8d", d => x"000dd7"),
    (y => x"a841ba", d => x"000dd3"),
    (y => x"a833e8", d => x"000dd2"),
    (y => x"a82618", d => x"000dd0"),
    (y => x"a8184b", d => x"000dcd"),
    (y => x"a80a81", d => x"000dca"),
    (y => x"a7fcb8", d => x"000dc9"),
    (y => x"a7eef2", d => x"000dc6"),
    (y => x"a7e12e", d => x"000dc4"),
    (y => x"a7d36c", d => x"000dc2"),
    (y => x"a7c5ac", d => x"000dc0"),
    (y => x"a7b7ef", d => x"000dbd"),
    (y => x"a7aa34", d => x"000dbb"),
    (y => x"a79c7b", d => x"000db9"),
    (y => x"a78ec4", d => x"000db7"),
    (y => x"a78110", d => x"000db4"),
    (y => x"a7735e", d => x"000db2"),
    (y => x"a765ae", d => x"000db0"),
    (y => x"a75801", d => x"000dad"),
    (y => x"a74a55", d => x"000dac"),
    (y => x"a73cac", d => x"000da9"),
    (y => x"a72f05", d => x"000da7"),
    (y => x"a72160", d => x"000da5"),
    (y => x"a713be", d => x"000da2"),
    (y => x"a7061e", d => x"000da0"),
    (y => x"a6f880", d => x"000d9e"),
    (y => x"a6eae4", d => x"000d9c"),
    (y => x"a6dd4a", d => x"000d9a"),
    (y => x"a6cfb3", d => x"000d97"),
    (y => x"a6c21e", d => x"000d95"),
    (y => x"a6b48b", d => x"000d93"),
    (y => x"a6a6fa", d => x"000d91"),
    (y => x"a6996c", d => x"000d8e"),
    (y => x"a68bdf", d => x"000d8d"),
    (y => x"a67e55", d => x"000d8a"),
    (y => x"a670cd", d => x"000d88"),
    (y => x"a66348", d => x"000d85"),
    (y => x"a655c4", d => x"000d84"),
    (y => x"a64843", d => x"000d81"),
    (y => x"a63ac4", d => x"000d7f"),
    (y => x"a62d47", d => x"000d7d"),
    (y => x"a61fcc", d => x"000d7b"),
    (y => x"a61253", d => x"000d79"),
    (y => x"a604dd", d => x"000d76"),
    (y => x"a5f769", d => x"000d74"),
    (y => x"a5e9f7", d => x"000d72"),
    (y => x"a5dc87", d => x"000d70"),
    (y => x"a5cf19", d => x"000d6e"),
    (y => x"a5c1ae", d => x"000d6b"),
    (y => x"a5b444", d => x"000d6a"),
    (y => x"a5a6dd", d => x"000d67"),
    (y => x"a59978", d => x"000d65"),
    (y => x"a58c16", d => x"000d62"),
    (y => x"a57eb5", d => x"000d61"),
    (y => x"a57156", d => x"000d5f"),
    (y => x"a563fa", d => x"000d5c"),
    (y => x"a556a0", d => x"000d5a"),
    (y => x"a54948", d => x"000d58"),
    (y => x"a53bf2", d => x"000d56"),
    (y => x"a52e9e", d => x"000d54"),
    (y => x"a5214d", d => x"000d51"),
    (y => x"a513fd", d => x"000d50"),
    (y => x"a506b0", d => x"000d4d"),
    (y => x"a4f965", d => x"000d4b"),
    (y => x"a4ec1c", d => x"000d49"),
    (y => x"a4ded5", d => x"000d47"),
    (y => x"a4d190", d => x"000d45"),
    (y => x"a4c44e", d => x"000d42"),
    (y => x"a4b70d", d => x"000d41"),
    (y => x"a4a9cf", d => x"000d3e"),
    (y => x"a49c93", d => x"000d3c"),
    (y => x"a48f59", d => x"000d3a"),
    (y => x"a48221", d => x"000d38"),
    (y => x"a474eb", d => x"000d36"),
    (y => x"a467b7", d => x"000d34"),
    (y => x"a45a86", d => x"000d31"),
    (y => x"a44d56", d => x"000d30"),
    (y => x"a44029", d => x"000d2d"),
    (y => x"a432fe", d => x"000d2b"),
    (y => x"a425d5", d => x"000d29"),
    (y => x"a418ae", d => x"000d27"),
    (y => x"a40b89", d => x"000d25"),
    (y => x"a3fe66", d => x"000d23"),
    (y => x"a3f145", d => x"000d21"),
    (y => x"a3e427", d => x"000d1e"),
    (y => x"a3d70a", d => x"000d1d"),
    (y => x"a3c9f0", d => x"000d1a"),
    (y => x"a3bcd7", d => x"000d19"),
    (y => x"a3afc1", d => x"000d16"),
    (y => x"a3a2ad", d => x"000d14"),
    (y => x"a3959b", d => x"000d12"),
    (y => x"a3888b", d => x"000d10"),
    (y => x"a37b7d", d => x"000d0e"),
    (y => x"a36e72", d => x"000d0b"),
    (y => x"a36168", d => x"000d0a"),
    (y => x"a35460", d => x"000d08"),
    (y => x"a3475b", d => x"000d05"),
    (y => x"a33a57", d => x"000d04"),
    (y => x"a32d56", d => x"000d01"),
    (y => x"a32057", d => x"000cff"),
    (y => x"a31359", d => x"000cfe"),
    (y => x"a3065e", d => x"000cfb"),
    (y => x"a2f965", d => x"000cf9"),
    (y => x"a2ec6e", d => x"000cf7"),
    (y => x"a2df79", d => x"000cf5"),
    (y => x"a2d286", d => x"000cf3"),
    (y => x"a2c595", d => x"000cf1"),
    (y => x"a2b8a6", d => x"000cef"),
    (y => x"a2abba", d => x"000cec"),
    (y => x"a29ecf", d => x"000ceb"),
    (y => x"a291e6", d => x"000ce9"),
    (y => x"a28500", d => x"000ce6"),
    (y => x"a2781b", d => x"000ce5"),
    (y => x"a26b39", d => x"000ce2"),
    (y => x"a25e58", d => x"000ce1"),
    (y => x"a2517a", d => x"000cde"),
    (y => x"a2449d", d => x"000cdd"),
    (y => x"a237c3", d => x"000cda"),
    (y => x"a22aeb", d => x"000cd8"),
    (y => x"a21e14", d => x"000cd7"),
    (y => x"a21140", d => x"000cd4"),
    (y => x"a2046e", d => x"000cd2"),
    (y => x"a1f79e", d => x"000cd0"),
    (y => x"a1ead0", d => x"000cce"),
    (y => x"a1de04", d => x"000ccc"),
    (y => x"a1d139", d => x"000ccb"),
    (y => x"a1c471", d => x"000cc8"),
    (y => x"a1b7ab", d => x"000cc6"),
    (y => x"a1aae7", d => x"000cc4"),
    (y => x"a19e25", d => x"000cc2"),
    (y => x"a19165", d => x"000cc0"),
    (y => x"a184a7", d => x"000cbe"),
    (y => x"a177eb", d => x"000cbc"),
    (y => x"a16b31", d => x"000cba"),
    (y => x"a15e79", d => x"000cb8"),
    (y => x"a151c3", d => x"000cb6"),
    (y => x"a1450f", d => x"000cb4"),
    (y => x"a1385d", d => x"000cb2"),
    (y => x"a12bad", d => x"000cb0"),
    (y => x"a11eff", d => x"000cae"),
    (y => x"a11253", d => x"000cac"),
    (y => x"a105a9", d => x"000caa"),
    (y => x"a0f901", d => x"000ca8"),
    (y => x"a0ec5b", d => x"000ca6"),
    (y => x"a0dfb7", d => x"000ca4"),
    (y => x"a0d315", d => x"000ca2"),
    (y => x"a0c675", d => x"000ca0"),
    (y => x"a0b9d7", d => x"000c9e"),
    (y => x"a0ad3b", d => x"000c9c"),
    (y => x"a0a0a1", d => x"000c9a"),
    (y => x"a09408", d => x"000c99"),
    (y => x"a08772", d => x"000c96"),
    (y => x"a07ade", d => x"000c94"),
    (y => x"a06e4c", d => x"000c92"),
    (y => x"a061bb", d => x"000c91"),
    (y => x"a0552d", d => x"000c8e"),
    (y => x"a048a1", d => x"000c8c"),
    (y => x"a03c16", d => x"000c8b"),
    (y => x"a02f8e", d => x"000c88"),
    (y => x"a02308", d => x"000c86"),
    (y => x"a01683", d => x"000c85"),
    (y => x"a00a01", d => x"000c82"),
    (y => x"9ffd80", d => x"000c81"),
    (y => x"9ff101", d => x"000c7f"),
    (y => x"9fe485", d => x"000c7c"),
    (y => x"9fd80a", d => x"000c7b"),
    (y => x"9fcb91", d => x"000c79"),
    (y => x"9fbf1a", d => x"000c77"),
    (y => x"9fb2a5", d => x"000c75"),
    (y => x"9fa632", d => x"000c73"),
    (y => x"9f99c1", d => x"000c71"),
    (y => x"9f8d52", d => x"000c6f"),
    (y => x"9f80e5", d => x"000c6d"),
    (y => x"9f747a", d => x"000c6b"),
    (y => x"9f6811", d => x"000c69"),
    (y => x"9f5ba9", d => x"000c68"),
    (y => x"9f4f44", d => x"000c65"),
    (y => x"9f42e0", d => x"000c64"),
    (y => x"9f367f", d => x"000c61"),
    (y => x"9f2a1f", d => x"000c60"),
    (y => x"9f1dc2", d => x"000c5d"),
    (y => x"9f1166", d => x"000c5c"),
    (y => x"9f050c", d => x"000c5a"),
    (y => x"9ef8b4", d => x"000c58"),
    (y => x"9eec5e", d => x"000c56"),
    (y => x"9ee00a", d => x"000c54"),
    (y => x"9ed3b8", d => x"000c52"),
    (y => x"9ec767", d => x"000c51"),
    (y => x"9ebb19", d => x"000c4e"),
    (y => x"9eaecc", d => x"000c4d"),
    (y => x"9ea282", d => x"000c4a"),
    (y => x"9e9639", d => x"000c49"),
    (y => x"9e89f2", d => x"000c47"),
    (y => x"9e7dae", d => x"000c44"),
    (y => x"9e716b", d => x"000c43"),
    (y => x"9e6529", d => x"000c42"),
    (y => x"9e58ea", d => x"000c3f"),
    (y => x"9e4cad", d => x"000c3d"),
    (y => x"9e4072", d => x"000c3b"),
    (y => x"9e3438", d => x"000c3a"),
    (y => x"9e2800", d => x"000c38"),
    (y => x"9e1bcb", d => x"000c35"),
    (y => x"9e0f97", d => x"000c34"),
    (y => x"9e0365", d => x"000c32"),
    (y => x"9df735", d => x"000c30"),
    (y => x"9deb07", d => x"000c2e"),
    (y => x"9ddeda", d => x"000c2d"),
    (y => x"9dd2b0", d => x"000c2a"),
    (y => x"9dc687", d => x"000c29"),
    (y => x"9dba61", d => x"000c26"),
    (y => x"9dae3c", d => x"000c25"),
    (y => x"9da219", d => x"000c23"),
    (y => x"9d95f8", d => x"000c21"),
    (y => x"9d89d8", d => x"000c20"),
    (y => x"9d7dbb", d => x"000c1d"),
    (y => x"9d71a0", d => x"000c1b"),
    (y => x"9d6586", d => x"000c1a"),
    (y => x"9d596e", d => x"000c18"),
    (y => x"9d4d58", d => x"000c16"),
    (y => x"9d4144", d => x"000c14"),
    (y => x"9d3532", d => x"000c12"),
    (y => x"9d2922", d => x"000c10"),
    (y => x"9d1d13", d => x"000c0f"),
    (y => x"9d1106", d => x"000c0d"),
    (y => x"9d04fc", d => x"000c0a"),
    (y => x"9cf8f3", d => x"000c09"),
    (y => x"9cecec", d => x"000c07"),
    (y => x"9ce0e6", d => x"000c06"),
    (y => x"9cd4e3", d => x"000c03"),
    (y => x"9cc8e1", d => x"000c02"),
    (y => x"9cbce2", d => x"000bff"),
    (y => x"9cb0e4", d => x"000bfe"),
    (y => x"9ca4e7", d => x"000bfd"),
    (y => x"9c98ed", d => x"000bfa"),
    (y => x"9c8cf5", d => x"000bf8"),
    (y => x"9c80fe", d => x"000bf7"),
    (y => x"9c7509", d => x"000bf5"),
    (y => x"9c6916", d => x"000bf3"),
    (y => x"9c5d25", d => x"000bf1"),
    (y => x"9c5136", d => x"000bef"),
    (y => x"9c4549", d => x"000bed"),
    (y => x"9c395d", d => x"000bec"),
    (y => x"9c2d73", d => x"000bea"),
    (y => x"9c218b", d => x"000be8"),
    (y => x"9c15a5", d => x"000be6"),
    (y => x"9c09c0", d => x"000be5"),
    (y => x"9bfdde", d => x"000be2"),
    (y => x"9bf1fd", d => x"000be1"),
    (y => x"9be61e", d => x"000bdf"),
    (y => x"9bda41", d => x"000bdd"),
    (y => x"9bce66", d => x"000bdb"),
    (y => x"9bc28c", d => x"000bda"),
    (y => x"9bb6b4", d => x"000bd8"),
    (y => x"9baade", d => x"000bd6"),
    (y => x"9b9f0a", d => x"000bd4"),
    (y => x"9b9338", d => x"000bd2"),
    (y => x"9b8767", d => x"000bd1"),
    (y => x"9b7b99", d => x"000bce"),
    (y => x"9b6fcc", d => x"000bcd"),
    (y => x"9b6400", d => x"000bcc"),
    (y => x"9b5837", d => x"000bc9"),
    (y => x"9b4c70", d => x"000bc7"),
    (y => x"9b40aa", d => x"000bc6"),
    (y => x"9b34e6", d => x"000bc4"),
    (y => x"9b2923", d => x"000bc3"),
    (y => x"9b1d63", d => x"000bc0"),
    (y => x"9b11a4", d => x"000bbf"),
    (y => x"9b05e7", d => x"000bbd"),
    (y => x"9afa2c", d => x"000bbb"),
    (y => x"9aee73", d => x"000bb9"),
    (y => x"9ae2bb", d => x"000bb8"),
    (y => x"9ad705", d => x"000bb6"),
    (y => x"9acb51", d => x"000bb4"),
    (y => x"9abf9f", d => x"000bb2"),
    (y => x"9ab3ef", d => x"000bb0"),
    (y => x"9aa840", d => x"000baf"),
    (y => x"9a9c93", d => x"000bad"),
    (y => x"9a90e8", d => x"000bab"),
    (y => x"9a853e", d => x"000baa"),
    (y => x"9a7997", d => x"000ba7"),
    (y => x"9a6df1", d => x"000ba6"),
    (y => x"9a624c", d => x"000ba5"),
    (y => x"9a56aa", d => x"000ba2"),
    (y => x"9a4b09", d => x"000ba1"),
    (y => x"9a3f6a", d => x"000b9f"),
    (y => x"9a33cd", d => x"000b9d"),
    (y => x"9a2832", d => x"000b9b"),
    (y => x"9a1c98", d => x"000b9a"),
    (y => x"9a1100", d => x"000b98"),
    (y => x"9a056a", d => x"000b96"),
    (y => x"99f9d6", d => x"000b94"),
    (y => x"99ee43", d => x"000b93"),
    (y => x"99e2b2", d => x"000b91"),
    (y => x"99d723", d => x"000b8f"),
    (y => x"99cb95", d => x"000b8e"),
    (y => x"99c00a", d => x"000b8b"),
    (y => x"99b47f", d => x"000b8b"),
    (y => x"99a8f7", d => x"000b88"),
    (y => x"999d71", d => x"000b86"),
    (y => x"9991ec", d => x"000b85"),
    (y => x"998669", d => x"000b83"),
    (y => x"997ae7", d => x"000b82"),
    (y => x"996f68", d => x"000b7f"),
    (y => x"9963ea", d => x"000b7e"),
    (y => x"99586e", d => x"000b7c"),
    (y => x"994cf3", d => x"000b7b"),
    (y => x"99417a", d => x"000b79"),
    (y => x"993603", d => x"000b77"),
    (y => x"992a8e", d => x"000b75"),
    (y => x"991f1a", d => x"000b74"),
    (y => x"9913a8", d => x"000b72"),
    (y => x"990838", d => x"000b70"),
    (y => x"98fcca", d => x"000b6e"),
    (y => x"98f15d", d => x"000b6d"),
    (y => x"98e5f2", d => x"000b6b"),
    (y => x"98da88", d => x"000b6a"),
    (y => x"98cf21", d => x"000b67"),
    (y => x"98c3bb", d => x"000b66"),
    (y => x"98b856", d => x"000b65"),
    (y => x"98acf4", d => x"000b62"),
    (y => x"98a193", d => x"000b61"),
    (y => x"989634", d => x"000b5f"),
    (y => x"988ad6", d => x"000b5e"),
    (y => x"987f7a", d => x"000b5c"),
    (y => x"987420", d => x"000b5a"),
    (y => x"9868c8", d => x"000b58"),
    (y => x"985d71", d => x"000b57"),
    (y => x"98521c", d => x"000b55"),
    (y => x"9846c9", d => x"000b53"),
    (y => x"983b77", d => x"000b52"),
    (y => x"983027", d => x"000b50"),
    (y => x"9824d9", d => x"000b4e"),
    (y => x"98198c", d => x"000b4d"),
    (y => x"980e41", d => x"000b4b"),
    (y => x"9802f8", d => x"000b49"),
    (y => x"97f7b0", d => x"000b48"),
    (y => x"97ec6a", d => x"000b46"),
    (y => x"97e126", d => x"000b44"),
    (y => x"97d5e4", d => x"000b42"),
    (y => x"97caa3", d => x"000b41"),
    (y => x"97bf63", d => x"000b40"),
    (y => x"97b426", d => x"000b3d"),
    (y => x"97a8ea", d => x"000b3c"),
    (y => x"979db0", d => x"000b3a"),
    (y => x"979277", d => x"000b39"),
    (y => x"978740", d => x"000b37"),
    (y => x"977c0b", d => x"000b35"),
    (y => x"9770d7", d => x"000b34"),
    (y => x"9765a5", d => x"000b32"),
    (y => x"975a75", d => x"000b30"),
    (y => x"974f46", d => x"000b2f"),
    (y => x"974419", d => x"000b2d"),
    (y => x"9738ee", d => x"000b2b"),
    (y => x"972dc4", d => x"000b2a"),
    (y => x"97229c", d => x"000b28"),
    (y => x"971776", d => x"000b26"),
    (y => x"970c51", d => x"000b25"),
    (y => x"97012e", d => x"000b23"),
    (y => x"96f60c", d => x"000b22"),
    (y => x"96eaed", d => x"000b1f"),
    (y => x"96dfce", d => x"000b1f"),
    (y => x"96d4b2", d => x"000b1c"),
    (y => x"96c997", d => x"000b1b"),
    (y => x"96be7e", d => x"000b19"),
    (y => x"96b366", d => x"000b18"),
    (y => x"96a850", d => x"000b16"),
    (y => x"969d3c", d => x"000b14"),
    (y => x"969229", d => x"000b13"),
    (y => x"968718", d => x"000b11"),
    (y => x"967c08", d => x"000b10"),
    (y => x"9670fa", d => x"000b0e"),
    (y => x"9665ee", d => x"000b0c"),
    (y => x"965ae3", d => x"000b0b"),
    (y => x"964fda", d => x"000b09"),
    (y => x"9644d3", d => x"000b07"),
    (y => x"9639cd", d => x"000b06"),
    (y => x"962ec9", d => x"000b04"),
    (y => x"9623c6", d => x"000b03"),
    (y => x"9618c5", d => x"000b01"),
    (y => x"960dc6", d => x"000aff"),
    (y => x"9602c8", d => x"000afe"),
    (y => x"95f7cc", d => x"000afc"),
    (y => x"95ecd2", d => x"000afa"),
    (y => x"95e1d9", d => x"000af9"),
    (y => x"95d6e2", d => x"000af7"),
    (y => x"95cbec", d => x"000af6"),
    (y => x"95c0f8", d => x"000af4"),
    (y => x"95b605", d => x"000af3"),
    (y => x"95ab15", d => x"000af0"),
    (y => x"95a025", d => x"000af0"),
    (y => x"959538", d => x"000aed"),
    (y => x"958a4c", d => x"000aec"),
    (y => x"957f61", d => x"000aeb"),
    (y => x"957478", d => x"000ae9"),
    (y => x"956991", d => x"000ae7"),
    (y => x"955eab", d => x"000ae6"),
    (y => x"9553c7", d => x"000ae4"),
    (y => x"9548e4", d => x"000ae3"),
    (y => x"953e04", d => x"000ae0"),
    (y => x"953324", d => x"000ae0"),
    (y => x"952846", d => x"000ade"),
    (y => x"951d6a", d => x"000adc"),
    (y => x"951290", d => x"000ada"),
    (y => x"9507b7", d => x"000ad9"),
    (y => x"94fcdf", d => x"000ad8"),
    (y => x"94f209", d => x"000ad6"),
    (y => x"94e735", d => x"000ad4"),
    (y => x"94dc62", d => x"000ad3"),
    (y => x"94d191", d => x"000ad1"),
    (y => x"94c6c1", d => x"000ad0"),
    (y => x"94bbf3", d => x"000ace"),
    (y => x"94b127", d => x"000acc"),
    (y => x"94a65c", d => x"000acb"),
    (y => x"949b93", d => x"000ac9"),
    (y => x"9490cb", d => x"000ac8"),
    (y => x"948605", d => x"000ac6"),
    (y => x"947b40", d => x"000ac5"),
    (y => x"94707d", d => x"000ac3"),
    (y => x"9465bc", d => x"000ac1"),
    (y => x"945afc", d => x"000ac0"),
    (y => x"94503d", d => x"000abf"),
    (y => x"944580", d => x"000abd"),
    (y => x"943ac5", d => x"000abb"),
    (y => x"94300b", d => x"000aba"),
    (y => x"942553", d => x"000ab8"),
    (y => x"941a9d", d => x"000ab6"),
    (y => x"940fe8", d => x"000ab5"),
    (y => x"940534", d => x"000ab4"),
    (y => x"93fa82", d => x"000ab2"),
    (y => x"93efd2", d => x"000ab0"),
    (y => x"93e523", d => x"000aaf"),
    (y => x"93da75", d => x"000aae"),
    (y => x"93cfca", d => x"000aab"),
    (y => x"93c51f", d => x"000aab"),
    (y => x"93ba77", d => x"000aa8"),
    (y => x"93afcf", d => x"000aa8"),
    (y => x"93a52a", d => x"000aa5"),
    (y => x"939a86", d => x"000aa4"),
    (y => x"938fe3", d => x"000aa3"),
    (y => x"938542", d => x"000aa1"),
    (y => x"937aa3", d => x"000a9f"),
    (y => x"937005", d => x"000a9e"),
    (y => x"936568", d => x"000a9d"),
    (y => x"935acd", d => x"000a9b"),
    (y => x"935034", d => x"000a99"),
    (y => x"93459c", d => x"000a98"),
    (y => x"933b05", d => x"000a97"),
    (y => x"933071", d => x"000a94"),
    (y => x"9325dd", d => x"000a94"),
    (y => x"931b4b", d => x"000a92"),
    (y => x"9310bb", d => x"000a90"),
    (y => x"93062c", d => x"000a8f"),
    (y => x"92fb9f", d => x"000a8d"),
    (y => x"92f113", d => x"000a8c"),
    (y => x"92e689", d => x"000a8a"),
    (y => x"92dc00", d => x"000a89"),
    (y => x"92d179", d => x"000a87"),
    (y => x"92c6f4", d => x"000a85"),
    (y => x"92bc6f", d => x"000a85"),
    (y => x"92b1ed", d => x"000a82"),
    (y => x"92a76c", d => x"000a81"),
    (y => x"929cec", d => x"000a80"),
    (y => x"92926e", d => x"000a7e"),
    (y => x"9287f1", d => x"000a7d"),
    (y => x"927d76", d => x"000a7b"),
    (y => x"9272fc", d => x"000a7a"),
    (y => x"926884", d => x"000a78"),
    (y => x"925e0d", d => x"000a77"),
    (y => x"925398", d => x"000a75"),
    (y => x"924924", d => x"000a74"),
    (y => x"923eb2", d => x"000a72"),
    (y => x"923442", d => x"000a70"),
    (y => x"9229d2", d => x"000a70"),
    (y => x"921f65", d => x"000a6d"),
    (y => x"9214f8", d => x"000a6d"),
    (y => x"920a8e", d => x"000a6a"),
    (y => x"920024", d => x"000a6a"),
    (y => x"91f5bd", d => x"000a67"),
    (y => x"91eb56", d => x"000a67"),
    (y => x"91e0f2", d => x"000a64"),
    (y => x"91d68e", d => x"000a64"),
    (y => x"91cc2c", d => x"000a62"),
    (y => x"91c1cc", d => x"000a60"),
    (y => x"91b76d", d => x"000a5f"),
    (y => x"91ad10", d => x"000a5d"),
    (y => x"91a2b4", d => x"000a5c"),
    (y => x"919859", d => x"000a5b"),
    (y => x"918e00", d => x"000a59"),
    (y => x"9183a9", d => x"000a57"),
    (y => x"917953", d => x"000a56"),
    (y => x"916efe", d => x"000a55"),
    (y => x"9164ab", d => x"000a53"),
    (y => x"915a59", d => x"000a52"),
    (y => x"915009", d => x"000a50"),
    (y => x"9145ba", d => x"000a4f"),
    (y => x"913b6d", d => x"000a4d"),
    (y => x"913121", d => x"000a4c"),
    (y => x"9126d7", d => x"000a4a"),
    (y => x"911c8e", d => x"000a49"),
    (y => x"911246", d => x"000a48"),
    (y => x"910800", d => x"000a46"),
    (y => x"90fdbc", d => x"000a44"),
    (y => x"90f379", d => x"000a43"),
    (y => x"90e937", d => x"000a42"),
    (y => x"90def7", d => x"000a40"),
    (y => x"90d4b8", d => x"000a3f"),
    (y => x"90ca7b", d => x"000a3d"),
    (y => x"90c03f", d => x"000a3c"),
    (y => x"90b605", d => x"000a3a"),
    (y => x"90abcc", d => x"000a39"),
    (y => x"90a194", d => x"000a38"),
    (y => x"90975e", d => x"000a36"),
    (y => x"908d2a", d => x"000a34"),
    (y => x"9082f7", d => x"000a33"),
    (y => x"9078c5", d => x"000a32"),
    (y => x"906e95", d => x"000a30"),
    (y => x"906466", d => x"000a2f"),
    (y => x"905a38", d => x"000a2e"),
    (y => x"90500c", d => x"000a2c"),
    (y => x"9045e2", d => x"000a2a"),
    (y => x"903bb9", d => x"000a29"),
    (y => x"903191", d => x"000a28"),
    (y => x"90276b", d => x"000a26"),
    (y => x"901d46", d => x"000a25"),
    (y => x"901322", d => x"000a24"),
    (y => x"900900", d => x"000a22"),
    (y => x"8ffee0", d => x"000a20"),
    (y => x"8ff4c1", d => x"000a1f"),
    (y => x"8feaa3", d => x"000a1e"),
    (y => x"8fe087", d => x"000a1c"),
    (y => x"8fd66c", d => x"000a1b"),
    (y => x"8fcc52", d => x"000a1a"),
    (y => x"8fc23a", d => x"000a18"),
    (y => x"8fb824", d => x"000a16"),
    (y => x"8fae0f", d => x"000a15"),
    (y => x"8fa3fb", d => x"000a14"),
    (y => x"8f99e8", d => x"000a13"),
    (y => x"8f8fd8", d => x"000a10"),
    (y => x"8f85c8", d => x"000a10"),
    (y => x"8f7bba", d => x"000a0e"),
    (y => x"8f71ad", d => x"000a0d"),
    (y => x"8f67a2", d => x"000a0b"),
    (y => x"8f5d98", d => x"000a0a"),
    (y => x"8f538f", d => x"000a09"),
    (y => x"8f4988", d => x"000a07"),
    (y => x"8f3f83", d => x"000a05"),
    (y => x"8f357e", d => x"000a05"),
    (y => x"8f2b7b", d => x"000a03"),
    (y => x"8f217a", d => x"000a01"),
    (y => x"8f177a", d => x"000a00"),
    (y => x"8f0d7b", d => x"0009ff"),
    (y => x"8f037e", d => x"0009fd"),
    (y => x"8ef982", d => x"0009fc"),
    (y => x"8eef87", d => x"0009fb"),
    (y => x"8ee58e", d => x"0009f9"),
    (y => x"8edb96", d => x"0009f8"),
    (y => x"8ed1a0", d => x"0009f6"),
    (y => x"8ec7ab", d => x"0009f5"),
    (y => x"8ebdb8", d => x"0009f3"),
    (y => x"8eb3c5", d => x"0009f3"),
    (y => x"8ea9d5", d => x"0009f0"),
    (y => x"8e9fe5", d => x"0009f0"),
    (y => x"8e95f7", d => x"0009ee"),
    (y => x"8e8c0a", d => x"0009ed"),
    (y => x"8e821f", d => x"0009eb"),
    (y => x"8e7835", d => x"0009ea"),
    (y => x"8e6e4d", d => x"0009e8"),
    (y => x"8e6466", d => x"0009e7"),
    (y => x"8e5a80", d => x"0009e6"),
    (y => x"8e509c", d => x"0009e4"),
    (y => x"8e46b9", d => x"0009e3"),
    (y => x"8e3cd7", d => x"0009e2"),
    (y => x"8e32f7", d => x"0009e0"),
    (y => x"8e2918", d => x"0009df"),
    (y => x"8e1f3a", d => x"0009de"),
    (y => x"8e155e", d => x"0009dc"),
    (y => x"8e0b83", d => x"0009db"),
    (y => x"8e01aa", d => x"0009d9"),
    (y => x"8df7d2", d => x"0009d8"),
    (y => x"8dedfb", d => x"0009d7"),
    (y => x"8de426", d => x"0009d5"),
    (y => x"8dda52", d => x"0009d4"),
    (y => x"8dd07f", d => x"0009d3"),
    (y => x"8dc6ae", d => x"0009d1"),
    (y => x"8dbcde", d => x"0009d0"),
    (y => x"8db310", d => x"0009ce"),
    (y => x"8da943", d => x"0009cd"),
    (y => x"8d9f77", d => x"0009cc"),
    (y => x"8d95ac", d => x"0009cb"),
    (y => x"8d8be3", d => x"0009c9"),
    (y => x"8d821b", d => x"0009c8"),
    (y => x"8d7855", d => x"0009c6"),
    (y => x"8d6e90", d => x"0009c5"),
    (y => x"8d64cc", d => x"0009c4"),
    (y => x"8d5b0a", d => x"0009c2"),
    (y => x"8d5149", d => x"0009c1"),
    (y => x"8d4789", d => x"0009c0"),
    (y => x"8d3dcb", d => x"0009be"),
    (y => x"8d340e", d => x"0009bd"),
    (y => x"8d2a52", d => x"0009bc"),
    (y => x"8d2098", d => x"0009ba"),
    (y => x"8d16df", d => x"0009b9"),
    (y => x"8d0d28", d => x"0009b7"),
    (y => x"8d0371", d => x"0009b7"),
    (y => x"8cf9bc", d => x"0009b5"),
    (y => x"8cf009", d => x"0009b3"),
    (y => x"8ce656", d => x"0009b3"),
    (y => x"8cdca6", d => x"0009b0"),
    (y => x"8cd2f6", d => x"0009b0"),
    (y => x"8cc948", d => x"0009ae"),
    (y => x"8cbf9b", d => x"0009ad"),
    (y => x"8cb5ef", d => x"0009ac"),
    (y => x"8cac45", d => x"0009aa"),
    (y => x"8ca29c", d => x"0009a9"),
    (y => x"8c98f4", d => x"0009a8"),
    (y => x"8c8f4e", d => x"0009a6"),
    (y => x"8c85a9", d => x"0009a5"),
    (y => x"8c7c05", d => x"0009a4"),
    (y => x"8c7263", d => x"0009a2"),
    (y => x"8c68c2", d => x"0009a1"),
    (y => x"8c5f22", d => x"0009a0"),
    (y => x"8c5584", d => x"00099e"),
    (y => x"8c4be7", d => x"00099d"),
    (y => x"8c424b", d => x"00099c"),
    (y => x"8c38b1", d => x"00099a"),
    (y => x"8c2f18", d => x"000999"),
    (y => x"8c2580", d => x"000998"),
    (y => x"8c1be9", d => x"000997"),
    (y => x"8c1254", d => x"000995"),
    (y => x"8c08c0", d => x"000994"),
    (y => x"8bff2e", d => x"000992"),
    (y => x"8bf59d", d => x"000991"),
    (y => x"8bec0d", d => x"000990"),
    (y => x"8be27e", d => x"00098f"),
    (y => x"8bd8f1", d => x"00098d"),
    (y => x"8bcf65", d => x"00098c"),
    (y => x"8bc5da", d => x"00098b"),
    (y => x"8bbc51", d => x"000989"),
    (y => x"8bb2c9", d => x"000988"),
    (y => x"8ba942", d => x"000987"),
    (y => x"8b9fbc", d => x"000986"),
    (y => x"8b9638", d => x"000984"),
    (y => x"8b8cb5", d => x"000983"),
    (y => x"8b8334", d => x"000981"),
    (y => x"8b79b3", d => x"000981"),
    (y => x"8b7034", d => x"00097f"),
    (y => x"8b66b6", d => x"00097e"),
    (y => x"8b5d3a", d => x"00097c"),
    (y => x"8b53bf", d => x"00097b"),
    (y => x"8b4a45", d => x"00097a"),
    (y => x"8b40cc", d => x"000979"),
    (y => x"8b3755", d => x"000977"),
    (y => x"8b2ddf", d => x"000976"),
    (y => x"8b246a", d => x"000975"),
    (y => x"8b1af7", d => x"000973"),
    (y => x"8b1185", d => x"000972"),
    (y => x"8b0814", d => x"000971"),
    (y => x"8afea4", d => x"000970"),
    (y => x"8af536", d => x"00096e"),
    (y => x"8aebc9", d => x"00096d"),
    (y => x"8ae25d", d => x"00096c"),
    (y => x"8ad8f3", d => x"00096a"),
    (y => x"8acf8a", d => x"000969"),
    (y => x"8ac622", d => x"000968"),
    (y => x"8abcbb", d => x"000967"),
    (y => x"8ab356", d => x"000965"),
    (y => x"8aa9f2", d => x"000964"),
    (y => x"8aa08f", d => x"000963"),
    (y => x"8a972d", d => x"000962"),
    (y => x"8a8dcd", d => x"000960"),
    (y => x"8a846e", d => x"00095f"),
    (y => x"8a7b10", d => x"00095e"),
    (y => x"8a71b4", d => x"00095c"),
    (y => x"8a6859", d => x"00095b"),
    (y => x"8a5eff", d => x"00095a"),
    (y => x"8a55a6", d => x"000959"),
    (y => x"8a4c4f", d => x"000957"),
    (y => x"8a42f8", d => x"000957"),
    (y => x"8a39a3", d => x"000955"),
    (y => x"8a3050", d => x"000953"),
    (y => x"8a26fd", d => x"000953"),
    (y => x"8a1dac", d => x"000951"),
    (y => x"8a145c", d => x"000950"),
    (y => x"8a0b0e", d => x"00094e"),
    (y => x"8a01c0", d => x"00094e"),
    (y => x"89f874", d => x"00094c"),
    (y => x"89ef29", d => x"00094b"),
    (y => x"89e5e0", d => x"000949"),
    (y => x"89dc98", d => x"000948"),
    (y => x"89d350", d => x"000948"),
    (y => x"89ca0b", d => x"000945"),
    (y => x"89c0c6", d => x"000945"),
    (y => x"89b783", d => x"000943"),
    (y => x"89ae40", d => x"000943"),
    (y => x"89a500", d => x"000940"),
    (y => x"899bc0", d => x"000940"),
    (y => x"899282", d => x"00093e"),
    (y => x"898944", d => x"00093e"),
    (y => x"898009", d => x"00093b"),
    (y => x"8976ce", d => x"00093b"),
    (y => x"896d94", d => x"00093a"),
    (y => x"89645c", d => x"000938"),
    (y => x"895b25", d => x"000937"),
    (y => x"8951f0", d => x"000935"),
    (y => x"8948bb", d => x"000935"),
    (y => x"893f88", d => x"000933"),
    (y => x"893656", d => x"000932"),
    (y => x"892d25", d => x"000931"),
    (y => x"8923f5", d => x"000930"),
    (y => x"891ac7", d => x"00092e"),
    (y => x"89119a", d => x"00092d"),
    (y => x"89086e", d => x"00092c"),
    (y => x"88ff44", d => x"00092a"),
    (y => x"88f61a", d => x"00092a"),
    (y => x"88ecf2", d => x"000928"),
    (y => x"88e3cb", d => x"000927"),
    (y => x"88daa5", d => x"000926"),
    (y => x"88d181", d => x"000924"),
    (y => x"88c85d", d => x"000924"),
    (y => x"88bf3b", d => x"000922"),
    (y => x"88b61a", d => x"000921"),
    (y => x"88acfb", d => x"00091f"),
    (y => x"88a3dc", d => x"00091f"),
    (y => x"889abf", d => x"00091d"),
    (y => x"8891a3", d => x"00091c"),
    (y => x"888888", d => x"00091b"),
    (y => x"887f6f", d => x"000919"),
    (y => x"887657", d => x"000918"),
    (y => x"886d3f", d => x"000918"),
    (y => x"886429", d => x"000916"),
    (y => x"885b15", d => x"000914"),
    (y => x"885201", d => x"000914"),
    (y => x"8848ef", d => x"000912"),
    (y => x"883fde", d => x"000911"),
    (y => x"8836ce", d => x"000910"),
    (y => x"882dbf", d => x"00090f"),
    (y => x"8824b2", d => x"00090d"),
    (y => x"881ba6", d => x"00090c"),
    (y => x"88129a", d => x"00090c"),
    (y => x"880991", d => x"000909"),
    (y => x"880088", d => x"000909"),
    (y => x"87f780", d => x"000908"),
    (y => x"87ee7a", d => x"000906"),
    (y => x"87e575", d => x"000905"),
    (y => x"87dc71", d => x"000904"),
    (y => x"87d36f", d => x"000902"),
    (y => x"87ca6d", d => x"000902"),
    (y => x"87c16d", d => x"000900"),
    (y => x"87b86e", d => x"0008ff"),
    (y => x"87af70", d => x"0008fe"),
    (y => x"87a673", d => x"0008fd"),
    (y => x"879d78", d => x"0008fb"),
    (y => x"87947d", d => x"0008fb"),
    (y => x"878b84", d => x"0008f9"),
    (y => x"87828c", d => x"0008f8"),
    (y => x"877995", d => x"0008f7"),
    (y => x"8770a0", d => x"0008f5"),
    (y => x"8767ab", d => x"0008f5"),
    (y => x"875eb8", d => x"0008f3"),
    (y => x"8755c6", d => x"0008f2"),
    (y => x"874cd5", d => x"0008f1"),
    (y => x"8743e6", d => x"0008ef"),
    (y => x"873af7", d => x"0008ef"),
    (y => x"87320a", d => x"0008ed"),
    (y => x"87291e", d => x"0008ec"),
    (y => x"872033", d => x"0008eb"),
    (y => x"871749", d => x"0008ea"),
    (y => x"870e60", d => x"0008e9"),
    (y => x"870579", d => x"0008e7"),
    (y => x"86fc93", d => x"0008e6"),
    (y => x"86f3ad", d => x"0008e6"),
    (y => x"86eaca", d => x"0008e3"),
    (y => x"86e1e7", d => x"0008e3"),
    (y => x"86d905", d => x"0008e2"),
    (y => x"86d025", d => x"0008e0"),
    (y => x"86c746", d => x"0008df"),
    (y => x"86be67", d => x"0008df"),
    (y => x"86b58b", d => x"0008dc"),
    (y => x"86acaf", d => x"0008dc"),
    (y => x"86a3d4", d => x"0008db"),
    (y => x"869afb", d => x"0008d9"),
    (y => x"869223", d => x"0008d8"),
    (y => x"86894c", d => x"0008d7"),
    (y => x"868076", d => x"0008d6"),
    (y => x"8677a1", d => x"0008d5"),
    (y => x"866ecd", d => x"0008d4"),
    (y => x"8665fb", d => x"0008d2"),
    (y => x"865d2a", d => x"0008d1"),
    (y => x"865459", d => x"0008d1"),
    (y => x"864b8a", d => x"0008cf"),
    (y => x"8642bd", d => x"0008cd"),
    (y => x"8639f0", d => x"0008cd"),
    (y => x"863124", d => x"0008cc"),
    (y => x"86285a", d => x"0008ca"),
    (y => x"861f91", d => x"0008c9"),
    (y => x"8616c9", d => x"0008c8"),
    (y => x"860e02", d => x"0008c7"),
    (y => x"86053c", d => x"0008c6"),
    (y => x"85fc78", d => x"0008c4"),
    (y => x"85f3b4", d => x"0008c4"),
    (y => x"85eaf2", d => x"0008c2"),
    (y => x"85e231", d => x"0008c1"),
    (y => x"85d971", d => x"0008c0"),
    (y => x"85d0b2", d => x"0008bf"),
    (y => x"85c7f4", d => x"0008be"),
    (y => x"85bf37", d => x"0008bd"),
    (y => x"85b67c", d => x"0008bb"),
    (y => x"85adc2", d => x"0008ba"),
    (y => x"85a508", d => x"0008ba"),
    (y => x"859c50", d => x"0008b8"),
    (y => x"859399", d => x"0008b7"),
    (y => x"858ae4", d => x"0008b5"),
    (y => x"85822f", d => x"0008b5"),
    (y => x"85797b", d => x"0008b4"),
    (y => x"8570c9", d => x"0008b2"),
    (y => x"856818", d => x"0008b1"),
    (y => x"855f68", d => x"0008b0"),
    (y => x"8556b9", d => x"0008af"),
    (y => x"854e0b", d => x"0008ae"),
    (y => x"85455e", d => x"0008ad"),
    (y => x"853cb3", d => x"0008ab"),
    (y => x"853408", d => x"0008ab"),
    (y => x"852b5f", d => x"0008a9"),
    (y => x"8522b7", d => x"0008a8"),
    (y => x"851a10", d => x"0008a7"),
    (y => x"85116a", d => x"0008a6"),
    (y => x"8508c5", d => x"0008a5"),
    (y => x"850021", d => x"0008a4"),
    (y => x"84f77f", d => x"0008a2"),
    (y => x"84eedd", d => x"0008a2"),
    (y => x"84e63d", d => x"0008a0"),
    (y => x"84dd9e", d => x"00089f"),
    (y => x"84d4ff", d => x"00089f"),
    (y => x"84cc62", d => x"00089d"),
    (y => x"84c3c7", d => x"00089b"),
    (y => x"84bb2c", d => x"00089b"),
    (y => x"84b292", d => x"00089a"),
    (y => x"84a9fa", d => x"000898"),
    (y => x"84a162", d => x"000898"),
    (y => x"8498cc", d => x"000896"),
    (y => x"849037", d => x"000895"),
    (y => x"8487a3", d => x"000894"),
    (y => x"847f10", d => x"000893"),
    (y => x"84767e", d => x"000892"),
    (y => x"846ded", d => x"000891"),
    (y => x"84655e", d => x"00088f"),
    (y => x"845ccf", d => x"00088f"),
    (y => x"845442", d => x"00088d"),
    (y => x"844bb5", d => x"00088d"),
    (y => x"84432a", d => x"00088b"),
    (y => x"843aa0", d => x"00088a"),
    (y => x"843217", d => x"000889"),
    (y => x"84298f", d => x"000888"),
    (y => x"842108", d => x"000887"),
    (y => x"841882", d => x"000886"),
    (y => x"840ffe", d => x"000884"),
    (y => x"84077a", d => x"000884"),
    (y => x"83fef8", d => x"000882"),
    (y => x"83f677", d => x"000881"),
    (y => x"83edf6", d => x"000881"),
    (y => x"83e577", d => x"00087f"),
    (y => x"83dcf9", d => x"00087e"),
    (y => x"83d47c", d => x"00087d"),
    (y => x"83cc00", d => x"00087c"),
    (y => x"83c386", d => x"00087a"),
    (y => x"83bb0c", d => x"00087a"),
    (y => x"83b293", d => x"000879"),
    (y => x"83aa1c", d => x"000877"),
    (y => x"83a1a6", d => x"000876"),
    (y => x"839930", d => x"000876"),
    (y => x"8390bc", d => x"000874"),
    (y => x"838849", d => x"000873"),
    (y => x"837fd7", d => x"000872"),
    (y => x"837766", d => x"000871"),
    (y => x"836ef6", d => x"000870"),
    (y => x"836687", d => x"00086f"),
    (y => x"835e19", d => x"00086e"),
    (y => x"8355ad", d => x"00086c"),
    (y => x"834d41", d => x"00086c"),
    (y => x"8344d7", d => x"00086a"),
    (y => x"833c6d", d => x"00086a"),
    (y => x"833405", d => x"000868"),
    (y => x"832b9e", d => x"000867"),
    (y => x"832338", d => x"000866"),
    (y => x"831ad3", d => x"000865"),
    (y => x"83126f", d => x"000864"),
    (y => x"830a0c", d => x"000863"),
    (y => x"8301aa", d => x"000862"),
    (y => x"82f949", d => x"000861"),
    (y => x"82f0e9", d => x"000860"),
    (y => x"82e88b", d => x"00085e"),
    (y => x"82e02d", d => x"00085e"),
    (y => x"82d7d0", d => x"00085d"),
    (y => x"82cf75", d => x"00085b"),
    (y => x"82c71b", d => x"00085a"),
    (y => x"82bec1", d => x"00085a"),
    (y => x"82b669", d => x"000858"),
    (y => x"82ae12", d => x"000857"),
    (y => x"82a5bc", d => x"000856"),
    (y => x"829d67", d => x"000855"),
    (y => x"829513", d => x"000854"),
    (y => x"828cc0", d => x"000853"),
    (y => x"82846e", d => x"000852"),
    (y => x"827c1d", d => x"000851"),
    (y => x"8273cd", d => x"000850"),
    (y => x"826b7f", d => x"00084e"),
    (y => x"826331", d => x"00084e"),
    (y => x"825ae4", d => x"00084d"),
    (y => x"825299", d => x"00084b"),
    (y => x"824a4e", d => x"00084b"),
    (y => x"824205", d => x"000849"),
    (y => x"8239bd", d => x"000848"),
    (y => x"823175", d => x"000848"),
    (y => x"82292f", d => x"000846"),
    (y => x"8220ea", d => x"000845"),
    (y => x"8218a6", d => x"000844"),
    (y => x"821062", d => x"000844"),
    (y => x"820820", d => x"000842"),
    (y => x"81ffdf", d => x"000841"),
    (y => x"81f79f", d => x"000840"),
    (y => x"81ef61", d => x"00083e"),
    (y => x"81e723", d => x"00083e"),
    (y => x"81dee6", d => x"00083d"),
    (y => x"81d6aa", d => x"00083c"),
    (y => x"81ce6f", d => x"00083b"),
    (y => x"81c636", d => x"000839"),
    (y => x"81bdfd", d => x"000839"),
    (y => x"81b5c5", d => x"000838"),
    (y => x"81ad8f", d => x"000836"),
    (y => x"81a559", d => x"000836"),
    (y => x"819d25", d => x"000834"),
    (y => x"8194f1", d => x"000834"),
    (y => x"818cbf", d => x"000832"),
    (y => x"81848e", d => x"000831"),
    (y => x"817c5d", d => x"000831"),
    (y => x"81742e", d => x"00082f"),
    (y => x"816c00", d => x"00082e"),
    (y => x"8163d2", d => x"00082e"),
    (y => x"815ba6", d => x"00082c"),
    (y => x"81537b", d => x"00082b"),
    (y => x"814b51", d => x"00082a"),
    (y => x"814328", d => x"000829"),
    (y => x"813b00", d => x"000828"),
    (y => x"8132d9", d => x"000827"),
    (y => x"812ab3", d => x"000826"),
    (y => x"81228e", d => x"000825"),
    (y => x"811a6a", d => x"000824"),
    (y => x"811247", d => x"000823"),
    (y => x"810a25", d => x"000822"),
    (y => x"810204", d => x"000821"),
    (y => x"80f9e4", d => x"000820"),
    (y => x"80f1c5", d => x"00081f"),
    (y => x"80e9a7", d => x"00081e"),
    (y => x"80e18b", d => x"00081c"),
    (y => x"80d96f", d => x"00081c"),
    (y => x"80d154", d => x"00081b"),
    (y => x"80c93a", d => x"00081a"),
    (y => x"80c122", d => x"000818"),
    (y => x"80b90a", d => x"000818"),
    (y => x"80b0f3", d => x"000817"),
    (y => x"80a8de", d => x"000815"),
    (y => x"80a0c9", d => x"000815"),
    (y => x"8098b5", d => x"000814"),
    (y => x"8090a3", d => x"000812"),
    (y => x"808891", d => x"000812"),
    (y => x"808080", d => x"000811"),
    (y => x"807871", d => x"00080f"),
    (y => x"807062", d => x"00080f"),
    (y => x"806855", d => x"00080d"),
    (y => x"806048", d => x"00080d"),
    (y => x"80583d", d => x"00080b"),
    (y => x"805032", d => x"00080b"),
    (y => x"804829", d => x"000809"),
    (y => x"804020", d => x"000809"),
    (y => x"803818", d => x"000808"),
    (y => x"803012", d => x"000806"),
    (y => x"80280c", d => x"000806"),
    (y => x"802008", d => x"000804"),
    (y => x"801804", d => x"000804"),
    (y => x"801002", d => x"000802"),
    (y => x"800800", d => x"000802"),
    (y => x"800000", d => x"000800"));

end package body;
