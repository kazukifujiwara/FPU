library IEEE;
use IEEE.std_logic_1164.all;

package finv_p is

  component finv is
    port (
      a : in std_logic_vector(31 downto 0);
      s : out std_logic_vector(31 downto 0));
  end component;

end package;


library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_misc.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

library work;
use work.fpu_util_p.all;

entity finv is
  port ( A : in  std_logic_vector(31 downto 0);
         S : out std_logic_vector(31 downto 0));
end entity finv;

architecture blackbox of FINV is

  -- a(32bit) & b(32bit) の計64bitを返す
  function table(index: std_logic_vector(10 downto 0))
    return std_logic_vector
  is
    variable r : std_logic_vector(63 downto 0);
  begin
    case conv_integer(index) is
      when    0 => r := x"3f7fe0043ffff002";
      when    1 => r := x"3f7fa01c3fffd00a";
      when    2 => r := x"3f7f604c3fffb01a";
      when    3 => r := x"3f7f20943fff9032";
      when    4 => r := x"3f7ee0f33fff7052";
      when    5 => r := x"3f7ea16b3fff5079";
      when    6 => r := x"3f7e61fa3fff30a9";
      when    7 => r := x"3f7e22a13fff10e1";
      when    8 => r := x"3f7de35f3ffef121";
      when    9 => r := x"3f7da4353ffed168";
      when   10 => r := x"3f7d65233ffeb1b7";
      when   11 => r := x"3f7d26283ffe920f";
      when   12 => r := x"3f7ce7453ffe726e";
      when   13 => r := x"3f7ca8793ffe52d5";
      when   14 => r := x"3f7c69c43ffe3344";
      when   15 => r := x"3f7c2b273ffe13bb";
      when   16 => r := x"3f7beca13ffdf439";
      when   17 => r := x"3f7bae333ffdd4bf";
      when   18 => r := x"3f7b6fdb3ffdb54d";
      when   19 => r := x"3f7b319b3ffd95e3";
      when   20 => r := x"3f7af3713ffd7681";
      when   21 => r := x"3f7ab55f3ffd5727";
      when   22 => r := x"3f7a77643ffd37d4";
      when   23 => r := x"3f7a39803ffd1889";
      when   24 => r := x"3f79fbb33ffcf945";
      when   25 => r := x"3f79bdfc3ffcda0a";
      when   26 => r := x"3f79805d3ffcbad6";
      when   27 => r := x"3f7942d43ffc9baa";
      when   28 => r := x"3f7905623ffc7c85";
      when   29 => r := x"3f78c8073ffc5d68";
      when   30 => r := x"3f788ac23ffc3e53";
      when   31 => r := x"3f784d943ffc1f46";
      when   32 => r := x"3f78107d3ffc0040";
      when   33 => r := x"3f77d37c3ffbe141";
      when   34 => r := x"3f7796923ffbc24b";
      when   35 => r := x"3f7759be3ffba35c";
      when   36 => r := x"3f771d003ffb8474";
      when   37 => r := x"3f76e0593ffb6595";
      when   38 => r := x"3f76a3c83ffb46bc";
      when   39 => r := x"3f76674e3ffb27ec";
      when   40 => r := x"3f762ae93ffb0922";
      when   41 => r := x"3f75ee9b3ffaea61";
      when   42 => r := x"3f75b2633ffacba7";
      when   43 => r := x"3f7576413ffaacf4";
      when   44 => r := x"3f753a363ffa8e49";
      when   45 => r := x"3f74fe403ffa6fa6";
      when   46 => r := x"3f74c2603ffa510a";
      when   47 => r := x"3f7486963ffa3275";
      when   48 => r := x"3f744ae23ffa13e8";
      when   49 => r := x"3f740f443ff9f562";
      when   50 => r := x"3f73d3bc3ff9d6e4";
      when   51 => r := x"3f7398493ff9b86d";
      when   52 => r := x"3f735ced3ff999fe";
      when   53 => r := x"3f7321a53ff97b96";
      when   54 => r := x"3f72e6743ff95d36";
      when   55 => r := x"3f72ab583ff93edd";
      when   56 => r := x"3f7270523ff9208b";
      when   57 => r := x"3f7235613ff90241";
      when   58 => r := x"3f71fa863ff8e3fe";
      when   59 => r := x"3f71bfc03ff8c5c2";
      when   60 => r := x"3f7185103ff8a78e";
      when   61 => r := x"3f714a743ff88961";
      when   62 => r := x"3f710fef3ff86b3b";
      when   63 => r := x"3f70d57e3ff84d1d";
      when   64 => r := x"3f709b233ff82f06";
      when   65 => r := x"3f7060dd3ff810f6";
      when   66 => r := x"3f7026ac3ff7f2ed";
      when   67 => r := x"3f6fec903ff7d4ec";
      when   68 => r := x"3f6fb28a3ff7b6f2";
      when   69 => r := x"3f6f78983ff79900";
      when   70 => r := x"3f6f3ebb3ff77b14";
      when   71 => r := x"3f6f04f43ff75d30";
      when   72 => r := x"3f6ecb413ff73f53";
      when   73 => r := x"3f6e91a33ff7217d";
      when   74 => r := x"3f6e581a3ff703ae";
      when   75 => r := x"3f6e1ea63ff6e5e7";
      when   76 => r := x"3f6de5473ff6c827";
      when   77 => r := x"3f6dabfc3ff6aa6e";
      when   78 => r := x"3f6d72c63ff68cbc";
      when   79 => r := x"3f6d39a43ff66f11";
      when   80 => r := x"3f6d00983ff6516d";
      when   81 => r := x"3f6cc79f3ff633d1";
      when   82 => r := x"3f6c8ebc3ff6163b";
      when   83 => r := x"3f6c55ed3ff5f8ad";
      when   84 => r := x"3f6c1d323ff5db26";
      when   85 => r := x"3f6be48b3ff5bda6";
      when   86 => r := x"3f6babfa3ff5a02d";
      when   87 => r := x"3f6b737c3ff582bb";
      when   88 => r := x"3f6b3b133ff56550";
      when   89 => r := x"3f6b02be3ff547ec";
      when   90 => r := x"3f6aca7d3ff52a8f";
      when   91 => r := x"3f6a92503ff50d39";
      when   92 => r := x"3f6a5a383ff4efeb";
      when   93 => r := x"3f6a22333ff4d2a3";
      when   94 => r := x"3f69ea433ff4b562";
      when   95 => r := x"3f69b2673ff49828";
      when   96 => r := x"3f697a9f3ff47af5";
      when   97 => r := x"3f6942ea3ff45dca";
      when   98 => r := x"3f690b4a3ff440a5";
      when   99 => r := x"3f68d3be3ff42387";
      when  100 => r := x"3f689c453ff40670";
      when  101 => r := x"3f6864e03ff3e960";
      when  102 => r := x"3f682d8f3ff3cc57";
      when  103 => r := x"3f67f6523ff3af54";
      when  104 => r := x"3f67bf283ff39259";
      when  105 => r := x"3f6788123ff37565";
      when  106 => r := x"3f6751103ff35877";
      when  107 => r := x"3f671a213ff33b90";
      when  108 => r := x"3f66e3463ff31eb0";
      when  109 => r := x"3f66ac7f3ff301d7";
      when  110 => r := x"3f6675cb3ff2e505";
      when  111 => r := x"3f663f2a3ff2c83a";
      when  112 => r := x"3f66089d3ff2ab76";
      when  113 => r := x"3f65d2233ff28eb8";
      when  114 => r := x"3f659bbc3ff27201";
      when  115 => r := x"3f6565693ff25551";
      when  116 => r := x"3f652f293ff238a8";
      when  117 => r := x"3f64f8fc3ff21c05";
      when  118 => r := x"3f64c2e33ff1ff69";
      when  119 => r := x"3f648cdc3ff1e2d4";
      when  120 => r := x"3f6456e93ff1c646";
      when  121 => r := x"3f6421093ff1a9bf";
      when  122 => r := x"3f63eb3c3ff18d3e";
      when  123 => r := x"3f63b5823ff170c4";
      when  124 => r := x"3f637fdb3ff15451";
      when  125 => r := x"3f634a473ff137e4";
      when  126 => r := x"3f6314c63ff11b7e";
      when  127 => r := x"3f62df573ff0ff1f";
      when  128 => r := x"3f62a9fc3ff0e2c6";
      when  129 => r := x"3f6274b33ff0c674";
      when  130 => r := x"3f623f7d3ff0aa29";
      when  131 => r := x"3f620a5a3ff08de4";
      when  132 => r := x"3f61d54a3ff071a6";
      when  133 => r := x"3f61a04c3ff0556f";
      when  134 => r := x"3f616b613ff0393e";
      when  135 => r := x"3f6136893ff01d14";
      when  136 => r := x"3f6101c33ff000f1";
      when  137 => r := x"3f60cd0f3fefe4d4";
      when  138 => r := x"3f60986f3fefc8bd";
      when  139 => r := x"3f6063e03fefacae";
      when  140 => r := x"3f602f643fef90a4";
      when  141 => r := x"3f5ffafb3fef74a2";
      when  142 => r := x"3f5fc6a43fef58a6";
      when  143 => r := x"3f5f925f3fef3cb0";
      when  144 => r := x"3f5f5e2c3fef20c1";
      when  145 => r := x"3f5f2a0c3fef04d9";
      when  146 => r := x"3f5ef5fe3feee8f7";
      when  147 => r := x"3f5ec2023feecd1b";
      when  148 => r := x"3f5e8e193feeb146";
      when  149 => r := x"3f5e5a413fee9577";
      when  150 => r := x"3f5e267c3fee79af";
      when  151 => r := x"3f5df2c83fee5dee";
      when  152 => r := x"3f5dbf273fee4233";
      when  153 => r := x"3f5d8b983fee267e";
      when  154 => r := x"3f5d581b3fee0ad0";
      when  155 => r := x"3f5d24af3fedef28";
      when  156 => r := x"3f5cf1563fedd387";
      when  157 => r := x"3f5cbe0e3fedb7ec";
      when  158 => r := x"3f5c8ad83fed9c57";
      when  159 => r := x"3f5c57b53fed80c9";
      when  160 => r := x"3f5c24a23fed6541";
      when  161 => r := x"3f5bf1a23fed49c0";
      when  162 => r := x"3f5bbeb33fed2e45";
      when  163 => r := x"3f5b8bd63fed12d0";
      when  164 => r := x"3f5b590b3fecf762";
      when  165 => r := x"3f5b26513fecdbfa";
      when  166 => r := x"3f5af3a93fecc098";
      when  167 => r := x"3f5ac1133feca53d";
      when  168 => r := x"3f5a8e8e3fec89e8";
      when  169 => r := x"3f5a5c1a3fec6e99";
      when  170 => r := x"3f5a29b83fec5351";
      when  171 => r := x"3f59f7673fec380f";
      when  172 => r := x"3f59c5283fec1cd3";
      when  173 => r := x"3f5992fa3fec019e";
      when  174 => r := x"3f5960de3febe66e";
      when  175 => r := x"3f592ed23febcb45";
      when  176 => r := x"3f58fcd83febb023";
      when  177 => r := x"3f58caf03feb9506";
      when  178 => r := x"3f5899183feb79f0";
      when  179 => r := x"3f5867523feb5ee0";
      when  180 => r := x"3f58359d3feb43d6";
      when  181 => r := x"3f5803f93feb28d2";
      when  182 => r := x"3f57d2663feb0dd5";
      when  183 => r := x"3f57a0e43feaf2de";
      when  184 => r := x"3f576f733fead7ed";
      when  185 => r := x"3f573e133feabd02";
      when  186 => r := x"3f570cc43feaa21d";
      when  187 => r := x"3f56db863fea873f";
      when  188 => r := x"3f56aa593fea6c66";
      when  189 => r := x"3f56793d3fea5194";
      when  190 => r := x"3f5648313fea36c8";
      when  191 => r := x"3f5617373fea1c02";
      when  192 => r := x"3f55e64d3fea0142";
      when  193 => r := x"3f55b5743fe9e689";
      when  194 => r := x"3f5584ac3fe9cbd5";
      when  195 => r := x"3f5553f43fe9b127";
      when  196 => r := x"3f55234d3fe99680";
      when  197 => r := x"3f54f2b73fe97bdf";
      when  198 => r := x"3f54c2313fe96143";
      when  199 => r := x"3f5491bc3fe946ae";
      when  200 => r := x"3f5461573fe92c1f";
      when  201 => r := x"3f5431033fe91196";
      when  202 => r := x"3f5400c03fe8f713";
      when  203 => r := x"3f53d08d3fe8dc96";
      when  204 => r := x"3f53a06a3fe8c21e";
      when  205 => r := x"3f5370583fe8a7ad";
      when  206 => r := x"3f5340563fe88d42";
      when  207 => r := x"3f5310643fe872dd";
      when  208 => r := x"3f52e0833fe8587e";
      when  209 => r := x"3f52b0b23fe83e25";
      when  210 => r := x"3f5280f13fe823d2";
      when  211 => r := x"3f5251413fe80985";
      when  212 => r := x"3f5221a13fe7ef3e";
      when  213 => r := x"3f51f2113fe7d4fd";
      when  214 => r := x"3f51c2913fe7bac1";
      when  215 => r := x"3f5193213fe7a08c";
      when  216 => r := x"3f5163c13fe7865c";
      when  217 => r := x"3f5134713fe76c33";
      when  218 => r := x"3f5105323fe7520f";
      when  219 => r := x"3f50d6023fe737f2";
      when  220 => r := x"3f50a6e23fe71dda";
      when  221 => r := x"3f5077d33fe703c8";
      when  222 => r := x"3f5048d33fe6e9bc";
      when  223 => r := x"3f5019e33fe6cfb6";
      when  224 => r := x"3f4feb033fe6b5b5";
      when  225 => r := x"3f4fbc323fe69bbb";
      when  226 => r := x"3f4f8d723fe681c6";
      when  227 => r := x"3f4f5ec13fe667d8";
      when  228 => r := x"3f4f30203fe64def";
      when  229 => r := x"3f4f018f3fe6340c";
      when  230 => r := x"3f4ed30d3fe61a2e";
      when  231 => r := x"3f4ea49c3fe60057";
      when  232 => r := x"3f4e76393fe5e685";
      when  233 => r := x"3f4e47e73fe5ccb9";
      when  234 => r := x"3f4e19a43fe5b2f3";
      when  235 => r := x"3f4deb703fe59933";
      when  236 => r := x"3f4dbd4c3fe57f78";
      when  237 => r := x"3f4d8f383fe565c3";
      when  238 => r := x"3f4d61333fe54c14";
      when  239 => r := x"3f4d333d3fe5326b";
      when  240 => r := x"3f4d05573fe518c8";
      when  241 => r := x"3f4cd7813fe4ff2a";
      when  242 => r := x"3f4ca9b93fe4e592";
      when  243 => r := x"3f4c7c013fe4cbff";
      when  244 => r := x"3f4c4e593fe4b273";
      when  245 => r := x"3f4c20bf3fe498ec";
      when  246 => r := x"3f4bf3353fe47f6b";
      when  247 => r := x"3f4bc5ba3fe465ef";
      when  248 => r := x"3f4b984e3fe44c79";
      when  249 => r := x"3f4b6af23fe43309";
      when  250 => r := x"3f4b3da43fe4199e";
      when  251 => r := x"3f4b10663fe4003a";
      when  252 => r := x"3f4ae3373fe3e6da";
      when  253 => r := x"3f4ab6173fe3cd81";
      when  254 => r := x"3f4a89063fe3b42d";
      when  255 => r := x"3f4a5c043fe39ade";
      when  256 => r := x"3f4a2f113fe38196";
      when  257 => r := x"3f4a022d3fe36853";
      when  258 => r := x"3f49d5583fe34f15";
      when  259 => r := x"3f49a8923fe335dd";
      when  260 => r := x"3f497bda3fe31cab";
      when  261 => r := x"3f494f323fe3037e";
      when  262 => r := x"3f4922983fe2ea57";
      when  263 => r := x"3f48f60e3fe2d136";
      when  264 => r := x"3f48c9923fe2b81a";
      when  265 => r := x"3f489d243fe29f03";
      when  266 => r := x"3f4870c63fe285f2";
      when  267 => r := x"3f4844763fe26ce7";
      when  268 => r := x"3f4818353fe253e1";
      when  269 => r := x"3f47ec033fe23ae1";
      when  270 => r := x"3f47bfdf3fe221e6";
      when  271 => r := x"3f4793ca3fe208f1";
      when  272 => r := x"3f4767c33fe1f001";
      when  273 => r := x"3f473bcb3fe1d717";
      when  274 => r := x"3f470fe23fe1be32";
      when  275 => r := x"3f46e4073fe1a553";
      when  276 => r := x"3f46b83a3fe18c79";
      when  277 => r := x"3f468c7c3fe173a5";
      when  278 => r := x"3f4660cd3fe15ad6";
      when  279 => r := x"3f46352b3fe1420d";
      when  280 => r := x"3f4609993fe12949";
      when  281 => r := x"3f45de143fe1108b";
      when  282 => r := x"3f45b29e3fe0f7d1";
      when  283 => r := x"3f4587363fe0df1e";
      when  284 => r := x"3f455bdd3fe0c670";
      when  285 => r := x"3f4530923fe0adc7";
      when  286 => r := x"3f4505553fe09524";
      when  287 => r := x"3f44da263fe07c86";
      when  288 => r := x"3f44af053fe063ed";
      when  289 => r := x"3f4483f33fe04b5a";
      when  290 => r := x"3f4458ef3fe032cc";
      when  291 => r := x"3f442df93fe01a44";
      when  292 => r := x"3f4403113fe001c1";
      when  293 => r := x"3f43d8373fdfe943";
      when  294 => r := x"3f43ad6b3fdfd0ca";
      when  295 => r := x"3f4382ad3fdfb857";
      when  296 => r := x"3f4357fd3fdf9fea";
      when  297 => r := x"3f432d5b3fdf8781";
      when  298 => r := x"3f4302c73fdf6f1e";
      when  299 => r := x"3f42d8413fdf56c1";
      when  300 => r := x"3f42adc93fdf3e68";
      when  301 => r := x"3f42835e3fdf2615";
      when  302 => r := x"3f4259023fdf0dc8";
      when  303 => r := x"3f422eb33fdef57f";
      when  304 => r := x"3f4204733fdedd3c";
      when  305 => r := x"3f41da403fdec4fe";
      when  306 => r := x"3f41b01a3fdeacc5";
      when  307 => r := x"3f4186033fde9492";
      when  308 => r := x"3f415bf93fde7c64";
      when  309 => r := x"3f4131fd3fde643b";
      when  310 => r := x"3f41080f3fde4c17";
      when  311 => r := x"3f40de2e3fde33f9";
      when  312 => r := x"3f40b45b3fde1be0";
      when  313 => r := x"3f408a953fde03cc";
      when  314 => r := x"3f4060dd3fddebbd";
      when  315 => r := x"3f4037333fddd3b4";
      when  316 => r := x"3f400d963fddbbaf";
      when  317 => r := x"3f3fe4073fdda3b0";
      when  318 => r := x"3f3fba853fdd8bb6";
      when  319 => r := x"3f3f91103fdd73c2";
      when  320 => r := x"3f3f67a93fdd5bd2";
      when  321 => r := x"3f3f3e503fdd43e8";
      when  322 => r := x"3f3f15033fdd2c02";
      when  323 => r := x"3f3eebc53fdd1422";
      when  324 => r := x"3f3ec2933fdcfc47";
      when  325 => r := x"3f3e996f3fdce472";
      when  326 => r := x"3f3e70583fdccca1";
      when  327 => r := x"3f3e474f3fdcb4d6";
      when  328 => r := x"3f3e1e523fdc9d0f";
      when  329 => r := x"3f3df5633fdc854e";
      when  330 => r := x"3f3dcc813fdc6d92";
      when  331 => r := x"3f3da3ad3fdc55db";
      when  332 => r := x"3f3d7ae53fdc3e29";
      when  333 => r := x"3f3d522b3fdc267c";
      when  334 => r := x"3f3d297e3fdc0ed4";
      when  335 => r := x"3f3d00de3fdbf732";
      when  336 => r := x"3f3cd84b3fdbdf94";
      when  337 => r := x"3f3cafc53fdbc7fc";
      when  338 => r := x"3f3c874c3fdbb068";
      when  339 => r := x"3f3c5ee03fdb98da";
      when  340 => r := x"3f3c36813fdb8151";
      when  341 => r := x"3f3c0e2f3fdb69cc";
      when  342 => r := x"3f3be5ea3fdb524d";
      when  343 => r := x"3f3bbdb23fdb3ad3";
      when  344 => r := x"3f3b95873fdb235e";
      when  345 => r := x"3f3b6d693fdb0bed";
      when  346 => r := x"3f3b45573fdaf482";
      when  347 => r := x"3f3b1d533fdadd1c";
      when  348 => r := x"3f3af55b3fdac5bb";
      when  349 => r := x"3f3acd703fdaae5f";
      when  350 => r := x"3f3aa5923fda9708";
      when  351 => r := x"3f3a7dc03fda7fb5";
      when  352 => r := x"3f3a55fc3fda6868";
      when  353 => r := x"3f3a2e443fda5120";
      when  354 => r := x"3f3a06983fda39dd";
      when  355 => r := x"3f39defa3fda229e";
      when  356 => r := x"3f39b7683fda0b65";
      when  357 => r := x"3f398fe33fd9f430";
      when  358 => r := x"3f39686a3fd9dd01";
      when  359 => r := x"3f3940fe3fd9c5d6";
      when  360 => r := x"3f39199e3fd9aeb1";
      when  361 => r := x"3f38f24b3fd99790";
      when  362 => r := x"3f38cb053fd98074";
      when  363 => r := x"3f38a3cb3fd9695d";
      when  364 => r := x"3f387c9d3fd9524b";
      when  365 => r := x"3f38557c3fd93b3e";
      when  366 => r := x"3f382e683fd92436";
      when  367 => r := x"3f3807603fd90d32";
      when  368 => r := x"3f37e0643fd8f634";
      when  369 => r := x"3f37b9753fd8df3a";
      when  370 => r := x"3f3792923fd8c845";
      when  371 => r := x"3f376bbb3fd8b156";
      when  372 => r := x"3f3744f13fd89a6b";
      when  373 => r := x"3f371e333fd88384";
      when  374 => r := x"3f36f7813fd86ca3";
      when  375 => r := x"3f36d0db3fd855c6";
      when  376 => r := x"3f36aa423fd83eef";
      when  377 => r := x"3f3683b53fd8281c";
      when  378 => r := x"3f365d343fd8114e";
      when  379 => r := x"3f3636c03fd7fa85";
      when  380 => r := x"3f3610573fd7e3c0";
      when  381 => r := x"3f35e9fb3fd7cd01";
      when  382 => r := x"3f35c3ab3fd7b646";
      when  383 => r := x"3f359d663fd79f90";
      when  384 => r := x"3f35772e3fd788de";
      when  385 => r := x"3f3551023fd77232";
      when  386 => r := x"3f352ae23fd75b8a";
      when  387 => r := x"3f3504ce3fd744e7";
      when  388 => r := x"3f34dec63fd72e49";
      when  389 => r := x"3f34b8cb3fd717af";
      when  390 => r := x"3f3492da3fd7011b";
      when  391 => r := x"3f346cf63fd6ea8b";
      when  392 => r := x"3f34471e3fd6d3ff";
      when  393 => r := x"3f3421523fd6bd79";
      when  394 => r := x"3f33fb923fd6a6f7";
      when  395 => r := x"3f33d5dd3fd6907a";
      when  396 => r := x"3f33b0353fd67a02";
      when  397 => r := x"3f338a983fd6638e";
      when  398 => r := x"3f3365073fd64d1f";
      when  399 => r := x"3f333f813fd636b5";
      when  400 => r := x"3f331a083fd6204f";
      when  401 => r := x"3f32f49a3fd609ee";
      when  402 => r := x"3f32cf383fd5f392";
      when  403 => r := x"3f32a9e23fd5dd3a";
      when  404 => r := x"3f3284973fd5c6e7";
      when  405 => r := x"3f325f593fd5b099";
      when  406 => r := x"3f323a253fd59a50";
      when  407 => r := x"3f3214fe3fd5840b";
      when  408 => r := x"3f31efe23fd56dca";
      when  409 => r := x"3f31cad13fd5578f";
      when  410 => r := x"3f31a5cc3fd54158";
      when  411 => r := x"3f3180d33fd52b25";
      when  412 => r := x"3f315be53fd514f7";
      when  413 => r := x"3f3137033fd4fece";
      when  414 => r := x"3f31122c3fd4e8aa";
      when  415 => r := x"3f30ed613fd4d28a";
      when  416 => r := x"3f30c8a13fd4bc6e";
      when  417 => r := x"3f30a3ed3fd4a658";
      when  418 => r := x"3f307f443fd49045";
      when  419 => r := x"3f305aa63fd47a38";
      when  420 => r := x"3f3036143fd4642f";
      when  421 => r := x"3f30118e3fd44e2a";
      when  422 => r := x"3f2fed123fd4382a";
      when  423 => r := x"3f2fc8a23fd4222f";
      when  424 => r := x"3f2fa43d3fd40c38";
      when  425 => r := x"3f2f7fe43fd3f646";
      when  426 => r := x"3f2f5b963fd3e058";
      when  427 => r := x"3f2f37533fd3ca6f";
      when  428 => r := x"3f2f131b3fd3b48a";
      when  429 => r := x"3f2eeeef3fd39eaa";
      when  430 => r := x"3f2ecacd3fd388cf";
      when  431 => r := x"3f2ea6b73fd372f7";
      when  432 => r := x"3f2e82ac3fd35d25";
      when  433 => r := x"3f2e5ead3fd34757";
      when  434 => r := x"3f2e3ab83fd3318d";
      when  435 => r := x"3f2e16cf3fd31bc8";
      when  436 => r := x"3f2df2f03fd30608";
      when  437 => r := x"3f2dcf1d3fd2f04b";
      when  438 => r := x"3f2dab553fd2da94";
      when  439 => r := x"3f2d87983fd2c4e1";
      when  440 => r := x"3f2d63e53fd2af32";
      when  441 => r := x"3f2d403e3fd29988";
      when  442 => r := x"3f2d1ca23fd283e2";
      when  443 => r := x"3f2cf9113fd26e40";
      when  444 => r := x"3f2cd58b3fd258a4";
      when  445 => r := x"3f2cb20f3fd2430b";
      when  446 => r := x"3f2c8e9f3fd22d77";
      when  447 => r := x"3f2c6b3a3fd217e7";
      when  448 => r := x"3f2c47df3fd2025c";
      when  449 => r := x"3f2c248f3fd1ecd5";
      when  450 => r := x"3f2c014a3fd1d753";
      when  451 => r := x"3f2bde103fd1c1d5";
      when  452 => r := x"3f2bbae13fd1ac5c";
      when  453 => r := x"3f2b97bd3fd196e6";
      when  454 => r := x"3f2b74a33fd18176";
      when  455 => r := x"3f2b51943fd16c09";
      when  456 => r := x"3f2b2e903fd156a1";
      when  457 => r := x"3f2b0b973fd1413e";
      when  458 => r := x"3f2ae8a83fd12bde";
      when  459 => r := x"3f2ac5c43fd11683";
      when  460 => r := x"3f2aa2eb3fd1012d";
      when  461 => r := x"3f2a801c3fd0ebdb";
      when  462 => r := x"3f2a5d583fd0d68d";
      when  463 => r := x"3f2a3a9f3fd0c143";
      when  464 => r := x"3f2a17f03fd0abfe";
      when  465 => r := x"3f29f54c3fd096bd";
      when  466 => r := x"3f29d2b33fd08181";
      when  467 => r := x"3f29b0243fd06c49";
      when  468 => r := x"3f298d9f3fd05715";
      when  469 => r := x"3f296b253fd041e5";
      when  470 => r := x"3f2948b63fd02cba";
      when  471 => r := x"3f2926513fd01793";
      when  472 => r := x"3f2903f73fd00270";
      when  473 => r := x"3f28e1a73fcfed52";
      when  474 => r := x"3f28bf613fcfd838";
      when  475 => r := x"3f289d263fcfc322";
      when  476 => r := x"3f287af53fcfae11";
      when  477 => r := x"3f2858cf3fcf9903";
      when  478 => r := x"3f2836b33fcf83fb";
      when  479 => r := x"3f2814a13fcf6ef6";
      when  480 => r := x"3f27f29a3fcf59f5";
      when  481 => r := x"3f27d09d3fcf44f9";
      when  482 => r := x"3f27aeab3fcf3001";
      when  483 => r := x"3f278cc23fcf1b0d";
      when  484 => r := x"3f276ae43fcf061e";
      when  485 => r := x"3f2749113fcef133";
      when  486 => r := x"3f2727473fcedc4c";
      when  487 => r := x"3f2705883fcec769";
      when  488 => r := x"3f26e3d33fceb28a";
      when  489 => r := x"3f26c2283fce9db0";
      when  490 => r := x"3f26a0873fce88da";
      when  491 => r := x"3f267ef13fce7408";
      when  492 => r := x"3f265d653fce5f3a";
      when  493 => r := x"3f263be23fce4a71";
      when  494 => r := x"3f261a6a3fce35ab";
      when  495 => r := x"3f25f8fc3fce20ea";
      when  496 => r := x"3f25d7993fce0c2d";
      when  497 => r := x"3f25b63f3fcdf774";
      when  498 => r := x"3f2594ef3fcde2bf";
      when  499 => r := x"3f2573a93fcdce0f";
      when  500 => r := x"3f25526e3fcdb962";
      when  501 => r := x"3f25313c3fcda4ba";
      when  502 => r := x"3f2510143fcd9016";
      when  503 => r := x"3f24eef73fcd7b76";
      when  504 => r := x"3f24cde33fcd66da";
      when  505 => r := x"3f24acd93fcd5243";
      when  506 => r := x"3f248bd93fcd3daf";
      when  507 => r := x"3f246ae33fcd2920";
      when  508 => r := x"3f2449f73fcd1494";
      when  509 => r := x"3f2429153fcd000d";
      when  510 => r := x"3f24083d3fcceb8a";
      when  511 => r := x"3f23e76e3fccd70b";
      when  512 => r := x"3f23c6aa3fccc290";
      when  513 => r := x"3f23a5ef3fccae19";
      when  514 => r := x"3f23853e3fcc99a7";
      when  515 => r := x"3f2364973fcc8538";
      when  516 => r := x"3f2343f93fcc70ce";
      when  517 => r := x"3f2323663fcc5c67";
      when  518 => r := x"3f2302dc3fcc4805";
      when  519 => r := x"3f22e25b3fcc33a6";
      when  520 => r := x"3f22c1e53fcc1f4c";
      when  521 => r := x"3f22a1783fcc0af6";
      when  522 => r := x"3f2281153fcbf6a4";
      when  523 => r := x"3f2260bc3fcbe256";
      when  524 => r := x"3f22406c3fcbce0c";
      when  525 => r := x"3f2220263fcbb9c6";
      when  526 => r := x"3f21ffe93fcba584";
      when  527 => r := x"3f21dfb73fcb9146";
      when  528 => r := x"3f21bf8d3fcb7d0c";
      when  529 => r := x"3f219f6e3fcb68d6";
      when  530 => r := x"3f217f583fcb54a4";
      when  531 => r := x"3f215f4b3fcb4076";
      when  532 => r := x"3f213f483fcb2c4c";
      when  533 => r := x"3f211f4e3fcb1826";
      when  534 => r := x"3f20ff5e3fcb0404";
      when  535 => r := x"3f20df783fcaefe6";
      when  536 => r := x"3f20bf9b3fcadbcc";
      when  537 => r := x"3f209fc73fcac7b6";
      when  538 => r := x"3f207ffd3fcab3a4";
      when  539 => r := x"3f20603c3fca9f96";
      when  540 => r := x"3f2040853fca8b8c";
      when  541 => r := x"3f2020d73fca7786";
      when  542 => r := x"3f2001333fca6384";
      when  543 => r := x"3f1fe1983fca4f86";
      when  544 => r := x"3f1fc2063fca3b8c";
      when  545 => r := x"3f1fa27e3fca2795";
      when  546 => r := x"3f1f82ff3fca13a3";
      when  547 => r := x"3f1f63893fc9ffb5";
      when  548 => r := x"3f1f441c3fc9ebca";
      when  549 => r := x"3f1f24b93fc9d7e4";
      when  550 => r := x"3f1f055f3fc9c401";
      when  551 => r := x"3f1ee60f3fc9b022";
      when  552 => r := x"3f1ec6c73fc99c47";
      when  553 => r := x"3f1ea7893fc98871";
      when  554 => r := x"3f1e88543fc9749e";
      when  555 => r := x"3f1e69293fc960ce";
      when  556 => r := x"3f1e4a063fc94d03";
      when  557 => r := x"3f1e2aed3fc9393c";
      when  558 => r := x"3f1e0bdd3fc92579";
      when  559 => r := x"3f1decd63fc911b9";
      when  560 => r := x"3f1dcdd83fc8fdfd";
      when  561 => r := x"3f1daee33fc8ea46";
      when  562 => r := x"3f1d8ff73fc8d692";
      when  563 => r := x"3f1d71153fc8c2e2";
      when  564 => r := x"3f1d523b3fc8af35";
      when  565 => r := x"3f1d336b3fc89b8d";
      when  566 => r := x"3f1d14a33fc887e8";
      when  567 => r := x"3f1cf5e53fc87448";
      when  568 => r := x"3f1cd72f3fc860ab";
      when  569 => r := x"3f1cb8833fc84d12";
      when  570 => r := x"3f1c99e03fc8397d";
      when  571 => r := x"3f1c7b453fc825ec";
      when  572 => r := x"3f1c5cb43fc8125e";
      when  573 => r := x"3f1c3e2c3fc7fed4";
      when  574 => r := x"3f1c1fac3fc7eb4e";
      when  575 => r := x"3f1c01363fc7d7cc";
      when  576 => r := x"3f1be2c83fc7c44e";
      when  577 => r := x"3f1bc4633fc7b0d4";
      when  578 => r := x"3f1ba6073fc79d5d";
      when  579 => r := x"3f1b87b43fc789ea";
      when  580 => r := x"3f1b696a3fc7767b";
      when  581 => r := x"3f1b4b293fc76310";
      when  582 => r := x"3f1b2cf03fc74fa8";
      when  583 => r := x"3f1b0ec13fc73c45";
      when  584 => r := x"3f1af09a3fc728e5";
      when  585 => r := x"3f1ad27c3fc71588";
      when  586 => r := x"3f1ab4673fc70230";
      when  587 => r := x"3f1a965a3fc6eedb";
      when  588 => r := x"3f1a78563fc6db8a";
      when  589 => r := x"3f1a5a5b3fc6c83d";
      when  590 => r := x"3f1a3c693fc6b4f4";
      when  591 => r := x"3f1a1e7f3fc6a1ae";
      when  592 => r := x"3f1a009f3fc68e6c";
      when  593 => r := x"3f19e2c63fc67b2e";
      when  594 => r := x"3f19c4f73fc667f4";
      when  595 => r := x"3f19a7303fc654bd";
      when  596 => r := x"3f1989723fc6418a";
      when  597 => r := x"3f196bbc3fc62e5a";
      when  598 => r := x"3f194e0f3fc61b2f";
      when  599 => r := x"3f19306b3fc60807";
      when  600 => r := x"3f1912cf3fc5f4e3";
      when  601 => r := x"3f18f53c3fc5e1c2";
      when  602 => r := x"3f18d7b13fc5cea5";
      when  603 => r := x"3f18ba2f3fc5bb8c";
      when  604 => r := x"3f189cb63fc5a877";
      when  605 => r := x"3f187f453fc59565";
      when  606 => r := x"3f1861dc3fc58257";
      when  607 => r := x"3f18447c3fc56f4d";
      when  608 => r := x"3f1827253fc55c46";
      when  609 => r := x"3f1809d63fc54943";
      when  610 => r := x"3f17ec8f3fc53643";
      when  611 => r := x"3f17cf513fc52348";
      when  612 => r := x"3f17b21b3fc51050";
      when  613 => r := x"3f1794ee3fc4fd5b";
      when  614 => r := x"3f1777c93fc4ea6a";
      when  615 => r := x"3f175aad3fc4d77d";
      when  616 => r := x"3f173d993fc4c494";
      when  617 => r := x"3f17208d3fc4b1ae";
      when  618 => r := x"3f17038a3fc49ecc";
      when  619 => r := x"3f16e68f3fc48bed";
      when  620 => r := x"3f16c99d3fc47912";
      when  621 => r := x"3f16acb23fc4663b";
      when  622 => r := x"3f168fd03fc45367";
      when  623 => r := x"3f1672f73fc44097";
      when  624 => r := x"3f1656253fc42dca";
      when  625 => r := x"3f16395c3fc41b01";
      when  626 => r := x"3f161c9b3fc4083c";
      when  627 => r := x"3f15ffe33fc3f57a";
      when  628 => r := x"3f15e3333fc3e2bc";
      when  629 => r := x"3f15c68b3fc3d001";
      when  630 => r := x"3f15a9eb3fc3bd4a";
      when  631 => r := x"3f158d533fc3aa97";
      when  632 => r := x"3f1570c33fc397e7";
      when  633 => r := x"3f15543c3fc3853a";
      when  634 => r := x"3f1537bd3fc37292";
      when  635 => r := x"3f151b463fc35fec";
      when  636 => r := x"3f14fed73fc34d4b";
      when  637 => r := x"3f14e2703fc33aad";
      when  638 => r := x"3f14c6123fc32812";
      when  639 => r := x"3f14a9bb3fc3157b";
      when  640 => r := x"3f148d6d3fc302e8";
      when  641 => r := x"3f1471273fc2f058";
      when  642 => r := x"3f1454e83fc2ddcc";
      when  643 => r := x"3f1438b23fc2cb43";
      when  644 => r := x"3f141c843fc2b8bd";
      when  645 => r := x"3f14005e3fc2a63c";
      when  646 => r := x"3f13e4403fc293bd";
      when  647 => r := x"3f13c82a3fc28142";
      when  648 => r := x"3f13ac1c3fc26ecb";
      when  649 => r := x"3f1390163fc25c57";
      when  650 => r := x"3f1374183fc249e7";
      when  651 => r := x"3f1358213fc2377a";
      when  652 => r := x"3f133c333fc22511";
      when  653 => r := x"3f13204d3fc212ab";
      when  654 => r := x"3f13046f3fc20049";
      when  655 => r := x"3f12e8983fc1edea";
      when  656 => r := x"3f12ccca3fc1db8f";
      when  657 => r := x"3f12b1033fc1c937";
      when  658 => r := x"3f1295443fc1b6e3";
      when  659 => r := x"3f12798d3fc1a492";
      when  660 => r := x"3f125dde3fc19244";
      when  661 => r := x"3f1242373fc17ffa";
      when  662 => r := x"3f1226983fc16db4";
      when  663 => r := x"3f120b003fc15b71";
      when  664 => r := x"3f11ef713fc14931";
      when  665 => r := x"3f11d3e93fc136f5";
      when  666 => r := x"3f11b8693fc124bc";
      when  667 => r := x"3f119cf03fc11287";
      when  668 => r := x"3f1181803fc10055";
      when  669 => r := x"3f1166173fc0ee26";
      when  670 => r := x"3f114ab63fc0dbfb";
      when  671 => r := x"3f112f5c3fc0c9d4";
      when  672 => r := x"3f11140b3fc0b7af";
      when  673 => r := x"3f10f8c13fc0a58f";
      when  674 => r := x"3f10dd7f3fc09371";
      when  675 => r := x"3f10c2443fc08157";
      when  676 => r := x"3f10a7113fc06f41";
      when  677 => r := x"3f108be63fc05d2d";
      when  678 => r := x"3f1070c23fc04b1e";
      when  679 => r := x"3f1055a63fc03911";
      when  680 => r := x"3f103a923fc02708";
      when  681 => r := x"3f101f853fc01503";
      when  682 => r := x"3f1004803fc00300";
      when  683 => r := x"3f0fe9833fbff101";
      when  684 => r := x"3f0fce8d3fbfdf06";
      when  685 => r := x"3f0fb39f3fbfcd0e";
      when  686 => r := x"3f0f98b83fbfbb19";
      when  687 => r := x"3f0f7dd93fbfa928";
      when  688 => r := x"3f0f63013fbf973a";
      when  689 => r := x"3f0f48313fbf854f";
      when  690 => r := x"3f0f2d683fbf7368";
      when  691 => r := x"3f0f12a73fbf6184";
      when  692 => r := x"3f0ef7ee3fbf4fa3";
      when  693 => r := x"3f0edd3c3fbf3dc6";
      when  694 => r := x"3f0ec2913fbf2bec";
      when  695 => r := x"3f0ea7ee3fbf1a15";
      when  696 => r := x"3f0e8d523fbf0842";
      when  697 => r := x"3f0e72be3fbef672";
      when  698 => r := x"3f0e58313fbee4a5";
      when  699 => r := x"3f0e3dab3fbed2dc";
      when  700 => r := x"3f0e232d3fbec116";
      when  701 => r := x"3f0e08b73fbeaf53";
      when  702 => r := x"3f0dee483fbe9d93";
      when  703 => r := x"3f0dd3e03fbe8bd7";
      when  704 => r := x"3f0db97f3fbe7a1e";
      when  705 => r := x"3f0d9f263fbe6869";
      when  706 => r := x"3f0d84d43fbe56b7";
      when  707 => r := x"3f0d6a8a3fbe4508";
      when  708 => r := x"3f0d50473fbe335c";
      when  709 => r := x"3f0d360b3fbe21b4";
      when  710 => r := x"3f0d1bd63fbe100e";
      when  711 => r := x"3f0d01a93fbdfe6d";
      when  712 => r := x"3f0ce7833fbdecce";
      when  713 => r := x"3f0ccd643fbddb33";
      when  714 => r := x"3f0cb34d3fbdc99b";
      when  715 => r := x"3f0c993d3fbdb806";
      when  716 => r := x"3f0c7f343fbda674";
      when  717 => r := x"3f0c65323fbd94e6";
      when  718 => r := x"3f0c4b383fbd835b";
      when  719 => r := x"3f0c31443fbd71d3";
      when  720 => r := x"3f0c17583fbd604f";
      when  721 => r := x"3f0bfd733fbd4ecd";
      when  722 => r := x"3f0be3963fbd3d4f";
      when  723 => r := x"3f0bc9bf3fbd2bd5";
      when  724 => r := x"3f0baff03fbd1a5d";
      when  725 => r := x"3f0b96283fbd08e9";
      when  726 => r := x"3f0b7c663fbcf777";
      when  727 => r := x"3f0b62ac3fbce609";
      when  728 => r := x"3f0b48fa3fbcd49f";
      when  729 => r := x"3f0b2f4e3fbcc337";
      when  730 => r := x"3f0b15a93fbcb1d3";
      when  731 => r := x"3f0afc0c3fbca072";
      when  732 => r := x"3f0ae2753fbc8f14";
      when  733 => r := x"3f0ac8e63fbc7db9";
      when  734 => r := x"3f0aaf5d3fbc6c62";
      when  735 => r := x"3f0a95dc3fbc5b0d";
      when  736 => r := x"3f0a7c613fbc49bc";
      when  737 => r := x"3f0a62ee3fbc386e";
      when  738 => r := x"3f0a49823fbc2723";
      when  739 => r := x"3f0a301d3fbc15dc";
      when  740 => r := x"3f0a16be3fbc0497";
      when  741 => r := x"3f09fd673fbbf356";
      when  742 => r := x"3f09e4173fbbe218";
      when  743 => r := x"3f09cacd3fbbd0dd";
      when  744 => r := x"3f09b18b3fbbbfa5";
      when  745 => r := x"3f09984f3fbbae71";
      when  746 => r := x"3f097f1b3fbb9d3f";
      when  747 => r := x"3f0965ed3fbb8c11";
      when  748 => r := x"3f094cc73fbb7ae6";
      when  749 => r := x"3f0933a73fbb69be";
      when  750 => r := x"3f091a8e3fbb5899";
      when  751 => r := x"3f09017c3fbb4777";
      when  752 => r := x"3f08e8713fbb3659";
      when  753 => r := x"3f08cf6c3fbb253d";
      when  754 => r := x"3f08b66f3fbb1425";
      when  755 => r := x"3f089d783fbb030f";
      when  756 => r := x"3f0884893fbaf1fd";
      when  757 => r := x"3f086ba03fbae0ee";
      when  758 => r := x"3f0852be3fbacfe2";
      when  759 => r := x"3f0839e23fbabeda";
      when  760 => r := x"3f08210e3fbaadd4";
      when  761 => r := x"3f0808403fba9cd1";
      when  762 => r := x"3f07ef793fba8bd2";
      when  763 => r := x"3f07d6b93fba7ad5";
      when  764 => r := x"3f07be003fba69dc";
      when  765 => r := x"3f07a54d3fba58e6";
      when  766 => r := x"3f078ca13fba47f3";
      when  767 => r := x"3f0773fc3fba3703";
      when  768 => r := x"3f075b5d3fba2616";
      when  769 => r := x"3f0742c53fba152c";
      when  770 => r := x"3f072a343fba0445";
      when  771 => r := x"3f0711aa3fb9f361";
      when  772 => r := x"3f06f9263fb9e281";
      when  773 => r := x"3f06e0a93fb9d1a3";
      when  774 => r := x"3f06c8333fb9c0c9";
      when  775 => r := x"3f06afc33fb9aff1";
      when  776 => r := x"3f06975a3fb99f1d";
      when  777 => r := x"3f067ef83fb98e4b";
      when  778 => r := x"3f06669c3fb97d7d";
      when  779 => r := x"3f064e473fb96cb2";
      when  780 => r := x"3f0635f83fb95be9";
      when  781 => r := x"3f061db03fb94b24";
      when  782 => r := x"3f06056f3fb93a62";
      when  783 => r := x"3f05ed343fb929a3";
      when  784 => r := x"3f05d5003fb918e7";
      when  785 => r := x"3f05bcd23fb9082d";
      when  786 => r := x"3f05a4ab3fb8f777";
      when  787 => r := x"3f058c8a3fb8e6c4";
      when  788 => r := x"3f0574703fb8d614";
      when  789 => r := x"3f055c5c3fb8c567";
      when  790 => r := x"3f05444f3fb8b4bd";
      when  791 => r := x"3f052c493fb8a416";
      when  792 => r := x"3f0514493fb89372";
      when  793 => r := x"3f04fc4f3fb882d1";
      when  794 => r := x"3f04e45c3fb87233";
      when  795 => r := x"3f04cc6f3fb86198";
      when  796 => r := x"3f04b4893fb85100";
      when  797 => r := x"3f049caa3fb8406b";
      when  798 => r := x"3f0484d03fb82fd9";
      when  799 => r := x"3f046cfd3fb81f4a";
      when  800 => r := x"3f0455313fb80ebd";
      when  801 => r := x"3f043d6b3fb7fe34";
      when  802 => r := x"3f0425ab3fb7edae";
      when  803 => r := x"3f040df23fb7dd2b";
      when  804 => r := x"3f03f63f3fb7ccab";
      when  805 => r := x"3f03de933fb7bc2d";
      when  806 => r := x"3f03c6ed3fb7abb3";
      when  807 => r := x"3f03af4d3fb79b3c";
      when  808 => r := x"3f0397b43fb78ac7";
      when  809 => r := x"3f0380213fb77a56";
      when  810 => r := x"3f0368943fb769e7";
      when  811 => r := x"3f03510e3fb7597c";
      when  812 => r := x"3f03398e3fb74913";
      when  813 => r := x"3f0322143fb738ad";
      when  814 => r := x"3f030aa03fb7284a";
      when  815 => r := x"3f02f3333fb717ea";
      when  816 => r := x"3f02dbcc3fb7078e";
      when  817 => r := x"3f02c46c3fb6f734";
      when  818 => r := x"3f02ad113fb6e6dc";
      when  819 => r := x"3f0295bd3fb6d688";
      when  820 => r := x"3f027e703fb6c637";
      when  821 => r := x"3f0267283fb6b5e9";
      when  822 => r := x"3f024fe73fb6a59d";
      when  823 => r := x"3f0238ab3fb69555";
      when  824 => r := x"3f0221763fb6850f";
      when  825 => r := x"3f020a483fb674cc";
      when  826 => r := x"3f01f31f3fb6648c";
      when  827 => r := x"3f01dbfd3fb65450";
      when  828 => r := x"3f01c4e03fb64415";
      when  829 => r := x"3f01adca3fb633de";
      when  830 => r := x"3f0196bb3fb623aa";
      when  831 => r := x"3f017fb13fb61379";
      when  832 => r := x"3f0168ad3fb6034a";
      when  833 => r := x"3f0151b03fb5f31e";
      when  834 => r := x"3f013ab83fb5e2f6";
      when  835 => r := x"3f0123c73fb5d2d0";
      when  836 => r := x"3f010cdc3fb5c2ad";
      when  837 => r := x"3f00f5f73fb5b28d";
      when  838 => r := x"3f00df183fb5a26f";
      when  839 => r := x"3f00c83f3fb59255";
      when  840 => r := x"3f00b16d3fb5823d";
      when  841 => r := x"3f009aa03fb57228";
      when  842 => r := x"3f0083d93fb56216";
      when  843 => r := x"3f006d193fb55207";
      when  844 => r := x"3f00565e3fb541fb";
      when  845 => r := x"3f003faa3fb531f2";
      when  846 => r := x"3f0028fb3fb521eb";
      when  847 => r := x"3f0012533fb511e8";
      when  848 => r := x"3efff7603fb501e7";
      when  849 => r := x"3effca273fb4f1e9";
      when  850 => r := x"3eff9cfa3fb4e1ed";
      when  851 => r := x"3eff6fd93fb4d1f5";
      when  852 => r := x"3eff42c43fb4c1ff";
      when  853 => r := x"3eff15bb3fb4b20d";
      when  854 => r := x"3efee8be3fb4a21d";
      when  855 => r := x"3efebbcd3fb49230";
      when  856 => r := x"3efe8ee73fb48245";
      when  857 => r := x"3efe620e3fb4725e";
      when  858 => r := x"3efe35403fb46279";
      when  859 => r := x"3efe087e3fb45297";
      when  860 => r := x"3efddbc83fb442b8";
      when  861 => r := x"3efdaf1e3fb432dc";
      when  862 => r := x"3efd827f3fb42302";
      when  863 => r := x"3efd55ec3fb4132b";
      when  864 => r := x"3efd29653fb40357";
      when  865 => r := x"3efcfcea3fb3f386";
      when  866 => r := x"3efcd07b3fb3e3b8";
      when  867 => r := x"3efca4173fb3d3ec";
      when  868 => r := x"3efc77bf3fb3c423";
      when  869 => r := x"3efc4b723fb3b45d";
      when  870 => r := x"3efc1f313fb3a49a";
      when  871 => r := x"3efbf2fc3fb394d9";
      when  872 => r := x"3efbc6d33fb3851b";
      when  873 => r := x"3efb9ab53fb37560";
      when  874 => r := x"3efb6ea33fb365a8";
      when  875 => r := x"3efb429c3fb355f3";
      when  876 => r := x"3efb16a13fb34640";
      when  877 => r := x"3efaeab13fb33690";
      when  878 => r := x"3efabecd3fb326e2";
      when  879 => r := x"3efa92f43fb31738";
      when  880 => r := x"3efa67273fb30790";
      when  881 => r := x"3efa3b653fb2f7eb";
      when  882 => r := x"3efa0faf3fb2e849";
      when  883 => r := x"3ef9e4043fb2d8a9";
      when  884 => r := x"3ef9b8653fb2c90c";
      when  885 => r := x"3ef98cd13fb2b972";
      when  886 => r := x"3ef961493fb2a9da";
      when  887 => r := x"3ef935cc3fb29a46";
      when  888 => r := x"3ef90a5a3fb28ab4";
      when  889 => r := x"3ef8def43fb27b24";
      when  890 => r := x"3ef8b3993fb26b98";
      when  891 => r := x"3ef888493fb25c0e";
      when  892 => r := x"3ef85d053fb24c87";
      when  893 => r := x"3ef831cb3fb23d02";
      when  894 => r := x"3ef8069e3fb22d81";
      when  895 => r := x"3ef7db7b3fb21e02";
      when  896 => r := x"3ef7b0643fb20e85";
      when  897 => r := x"3ef785583fb1ff0c";
      when  898 => r := x"3ef75a573fb1ef95";
      when  899 => r := x"3ef72f613fb1e020";
      when  900 => r := x"3ef704773fb1d0af";
      when  901 => r := x"3ef6d9983fb1c140";
      when  902 => r := x"3ef6aec33fb1b1d3";
      when  903 => r := x"3ef683fa3fb1a26a";
      when  904 => r := x"3ef6593d3fb19303";
      when  905 => r := x"3ef62e8a3fb1839f";
      when  906 => r := x"3ef603e23fb1743d";
      when  907 => r := x"3ef5d9463fb164de";
      when  908 => r := x"3ef5aeb43fb15582";
      when  909 => r := x"3ef5842e3fb14628";
      when  910 => r := x"3ef559b23fb136d1";
      when  911 => r := x"3ef52f423fb1277d";
      when  912 => r := x"3ef504dd3fb1182b";
      when  913 => r := x"3ef4da823fb108dd";
      when  914 => r := x"3ef4b0333fb0f990";
      when  915 => r := x"3ef485ee3fb0ea46";
      when  916 => r := x"3ef45bb53fb0daff";
      when  917 => r := x"3ef431863fb0cbbb";
      when  918 => r := x"3ef407633fb0bc79";
      when  919 => r := x"3ef3dd4a3fb0ad3a";
      when  920 => r := x"3ef3b33c3fb09dfe";
      when  921 => r := x"3ef389393fb08ec4";
      when  922 => r := x"3ef35f413fb07f8c";
      when  923 => r := x"3ef335543fb07058";
      when  924 => r := x"3ef30b713fb06126";
      when  925 => r := x"3ef2e19a3fb051f6";
      when  926 => r := x"3ef2b7cd3fb042ca";
      when  927 => r := x"3ef28e0b3fb0339f";
      when  928 => r := x"3ef264543fb02478";
      when  929 => r := x"3ef23aa73fb01553";
      when  930 => r := x"3ef211053fb00630";
      when  931 => r := x"3ef1e76e3faff711";
      when  932 => r := x"3ef1bde23fafe7f4";
      when  933 => r := x"3ef194603fafd8d9";
      when  934 => r := x"3ef16ae93fafc9c1";
      when  935 => r := x"3ef1417d3fafbaac";
      when  936 => r := x"3ef1181c3fafab99";
      when  937 => r := x"3ef0eec53faf9c89";
      when  938 => r := x"3ef0c5783faf8d7b";
      when  939 => r := x"3ef09c373faf7e70";
      when  940 => r := x"3ef073003faf6f67";
      when  941 => r := x"3ef049d33faf6062";
      when  942 => r := x"3ef020b13faf515e";
      when  943 => r := x"3eeff79a3faf425d";
      when  944 => r := x"3eefce8d3faf335f";
      when  945 => r := x"3eefa58b3faf2464";
      when  946 => r := x"3eef7c933faf156b";
      when  947 => r := x"3eef53a53faf0674";
      when  948 => r := x"3eef2ac33faef780";
      when  949 => r := x"3eef01ea3faee88f";
      when  950 => r := x"3eeed91c3faed9a0";
      when  951 => r := x"3eeeb0593faecab4";
      when  952 => r := x"3eee87a03faebbca";
      when  953 => r := x"3eee5ef13faeace3";
      when  954 => r := x"3eee364d3fae9dfe";
      when  955 => r := x"3eee0db33fae8f1c";
      when  956 => r := x"3eede5243fae803c";
      when  957 => r := x"3eedbc9f3fae715f";
      when  958 => r := x"3eed94243fae6285";
      when  959 => r := x"3eed6bb43fae53ad";
      when  960 => r := x"3eed434e3fae44d7";
      when  961 => r := x"3eed1af23fae3604";
      when  962 => r := x"3eecf2a13fae2734";
      when  963 => r := x"3eecca593fae1866";
      when  964 => r := x"3eeca21d3fae099b";
      when  965 => r := x"3eec79ea3fadfad2";
      when  966 => r := x"3eec51c23fadec0b";
      when  967 => r := x"3eec29a33faddd47";
      when  968 => r := x"3eec018f3fadce86";
      when  969 => r := x"3eebd9863fadbfc7";
      when  970 => r := x"3eebb1863fadb10b";
      when  971 => r := x"3eeb89913fada251";
      when  972 => r := x"3eeb61a53fad939a";
      when  973 => r := x"3eeb39c43fad84e5";
      when  974 => r := x"3eeb11ed3fad7632";
      when  975 => r := x"3eeaea203fad6783";
      when  976 => r := x"3eeac25e3fad58d5";
      when  977 => r := x"3eea9aa53fad4a2a";
      when  978 => r := x"3eea72f63fad3b82";
      when  979 => r := x"3eea4b523fad2cdc";
      when  980 => r := x"3eea23b83fad1e38";
      when  981 => r := x"3ee9fc273fad0f97";
      when  982 => r := x"3ee9d4a13fad00f9";
      when  983 => r := x"3ee9ad243facf25d";
      when  984 => r := x"3ee985b23face3c3";
      when  985 => r := x"3ee95e493facd52c";
      when  986 => r := x"3ee936eb3facc697";
      when  987 => r := x"3ee90f973facb805";
      when  988 => r := x"3ee8e84c3faca976";
      when  989 => r := x"3ee8c10b3fac9ae8";
      when  990 => r := x"3ee899d53fac8c5d";
      when  991 => r := x"3ee872a83fac7dd5";
      when  992 => r := x"3ee84b853fac6f4f";
      when  993 => r := x"3ee8246c3fac60cc";
      when  994 => r := x"3ee7fd5d3fac524b";
      when  995 => r := x"3ee7d6583fac43cc";
      when  996 => r := x"3ee7af5c3fac3550";
      when  997 => r := x"3ee7886b3fac26d6";
      when  998 => r := x"3ee761833fac185f";
      when  999 => r := x"3ee73aa53fac09ea";
      when 1000 => r := x"3ee713d13fabfb77";
      when 1001 => r := x"3ee6ed063fabed07";
      when 1002 => r := x"3ee6c6463fabde9a";
      when 1003 => r := x"3ee69f8f3fabd02f";
      when 1004 => r := x"3ee678e23fabc1c6";
      when 1005 => r := x"3ee6523e3fabb35f";
      when 1006 => r := x"3ee62ba43faba4fb";
      when 1007 => r := x"3ee605143fab969a";
      when 1008 => r := x"3ee5de8e3fab883b";
      when 1009 => r := x"3ee5b8113fab79de";
      when 1010 => r := x"3ee5919e3fab6b84";
      when 1011 => r := x"3ee56b353fab5d2c";
      when 1012 => r := x"3ee544d53fab4ed6";
      when 1013 => r := x"3ee51e7f3fab4083";
      when 1014 => r := x"3ee4f8333fab3233";
      when 1015 => r := x"3ee4d1f03fab23e4";
      when 1016 => r := x"3ee4abb73fab1598";
      when 1017 => r := x"3ee485873fab074f";
      when 1018 => r := x"3ee45f613faaf908";
      when 1019 => r := x"3ee439443faaeac3";
      when 1020 => r := x"3ee413313faadc81";
      when 1021 => r := x"3ee3ed283faace41";
      when 1022 => r := x"3ee3c7283faac003";
      when 1023 => r := x"3ee3a1313faab1c8";
      when 1024 => r := x"3ee37b443faaa38f";
      when 1025 => r := x"3ee355603faa9558";
      when 1026 => r := x"3ee32f863faa8724";
      when 1027 => r := x"3ee309b63faa78f2";
      when 1028 => r := x"3ee2e3ee3faa6ac3";
      when 1029 => r := x"3ee2be313faa5c96";
      when 1030 => r := x"3ee2987c3faa4e6b";
      when 1031 => r := x"3ee272d13faa4043";
      when 1032 => r := x"3ee24d303faa321d";
      when 1033 => r := x"3ee227983faa23f9";
      when 1034 => r := x"3ee202093faa15d8";
      when 1035 => r := x"3ee1dc833faa07b9";
      when 1036 => r := x"3ee1b7073fa9f99c";
      when 1037 => r := x"3ee191943fa9eb82";
      when 1038 => r := x"3ee16c2b3fa9dd6a";
      when 1039 => r := x"3ee146cb3fa9cf54";
      when 1040 => r := x"3ee121743fa9c141";
      when 1041 => r := x"3ee0fc263fa9b330";
      when 1042 => r := x"3ee0d6e23fa9a522";
      when 1043 => r := x"3ee0b1a73fa99715";
      when 1044 => r := x"3ee08c753fa9890b";
      when 1045 => r := x"3ee0674c3fa97b04";
      when 1046 => r := x"3ee0422d3fa96cff";
      when 1047 => r := x"3ee01d173fa95efc";
      when 1048 => r := x"3edff80a3fa950fb";
      when 1049 => r := x"3edfd3063fa942fd";
      when 1050 => r := x"3edfae0b3fa93501";
      when 1051 => r := x"3edf891a3fa92707";
      when 1052 => r := x"3edf64313fa9190f";
      when 1053 => r := x"3edf3f523fa90b1a";
      when 1054 => r := x"3edf1a7c3fa8fd27";
      when 1055 => r := x"3edef5af3fa8ef37";
      when 1056 => r := x"3eded0eb3fa8e149";
      when 1057 => r := x"3edeac313fa8d35d";
      when 1058 => r := x"3ede877f3fa8c573";
      when 1059 => r := x"3ede62d63fa8b78c";
      when 1060 => r := x"3ede3e373fa8a9a7";
      when 1061 => r := x"3ede19a03fa89bc4";
      when 1062 => r := x"3eddf5133fa88de4";
      when 1063 => r := x"3eddd08e3fa88005";
      when 1064 => r := x"3eddac133fa8722a";
      when 1065 => r := x"3edd87a03fa86450";
      when 1066 => r := x"3edd63373fa85679";
      when 1067 => r := x"3edd3ed63fa848a4";
      when 1068 => r := x"3edd1a7f3fa83ad1";
      when 1069 => r := x"3edcf6303fa82d00";
      when 1070 => r := x"3edcd1eb3fa81f32";
      when 1071 => r := x"3edcadae3fa81166";
      when 1072 => r := x"3edc897a3fa8039c";
      when 1073 => r := x"3edc654f3fa7f5d5";
      when 1074 => r := x"3edc412d3fa7e810";
      when 1075 => r := x"3edc1d143fa7da4d";
      when 1076 => r := x"3edbf9043fa7cc8c";
      when 1077 => r := x"3edbd4fd3fa7bece";
      when 1078 => r := x"3edbb0fe3fa7b111";
      when 1079 => r := x"3edb8d083fa7a357";
      when 1080 => r := x"3edb691c3fa795a0";
      when 1081 => r := x"3edb45373fa787ea";
      when 1082 => r := x"3edb215c3fa77a37";
      when 1083 => r := x"3edafd8a3fa76c86";
      when 1084 => r := x"3edad9c03fa75ed7";
      when 1085 => r := x"3edab5ff3fa7512b";
      when 1086 => r := x"3eda92473fa74381";
      when 1087 => r := x"3eda6e983fa735d9";
      when 1088 => r := x"3eda4af13fa72833";
      when 1089 => r := x"3eda27533fa71a8f";
      when 1090 => r := x"3eda03be3fa70cee";
      when 1091 => r := x"3ed9e0313fa6ff4f";
      when 1092 => r := x"3ed9bcae3fa6f1b2";
      when 1093 => r := x"3ed999323fa6e417";
      when 1094 => r := x"3ed975c03fa6d67f";
      when 1095 => r := x"3ed952563fa6c8e8";
      when 1096 => r := x"3ed92ef53fa6bb54";
      when 1097 => r := x"3ed90b9c3fa6adc3";
      when 1098 => r := x"3ed8e84d3fa6a033";
      when 1099 => r := x"3ed8c5053fa692a6";
      when 1100 => r := x"3ed8a1c73fa6851a";
      when 1101 => r := x"3ed87e903fa67791";
      when 1102 => r := x"3ed85b633fa66a0b";
      when 1103 => r := x"3ed8383e3fa65c86";
      when 1104 => r := x"3ed815223fa64f03";
      when 1105 => r := x"3ed7f20e3fa64183";
      when 1106 => r := x"3ed7cf033fa63405";
      when 1107 => r := x"3ed7ac003fa62689";
      when 1108 => r := x"3ed789063fa61910";
      when 1109 => r := x"3ed766143fa60b98";
      when 1110 => r := x"3ed7432b3fa5fe23";
      when 1111 => r := x"3ed7204a3fa5f0b0";
      when 1112 => r := x"3ed6fd723fa5e33f";
      when 1113 => r := x"3ed6daa23fa5d5d0";
      when 1114 => r := x"3ed6b7da3fa5c864";
      when 1115 => r := x"3ed6951b3fa5baf9";
      when 1116 => r := x"3ed672653fa5ad91";
      when 1117 => r := x"3ed64fb73fa5a02b";
      when 1118 => r := x"3ed62d113fa592c7";
      when 1119 => r := x"3ed60a743fa58565";
      when 1120 => r := x"3ed5e7df3fa57806";
      when 1121 => r := x"3ed5c5533fa56aa8";
      when 1122 => r := x"3ed5a2ce3fa55d4d";
      when 1123 => r := x"3ed580533fa54ff4";
      when 1124 => r := x"3ed55ddf3fa5429d";
      when 1125 => r := x"3ed53b743fa53548";
      when 1126 => r := x"3ed519113fa527f6";
      when 1127 => r := x"3ed4f6b73fa51aa5";
      when 1128 => r := x"3ed4d4653fa50d57";
      when 1129 => r := x"3ed4b21b3fa5000b";
      when 1130 => r := x"3ed48fd93fa4f2c0";
      when 1131 => r := x"3ed46da03fa4e579";
      when 1132 => r := x"3ed44b6f3fa4d833";
      when 1133 => r := x"3ed429463fa4caef";
      when 1134 => r := x"3ed407263fa4bdae";
      when 1135 => r := x"3ed3e50d3fa4b06e";
      when 1136 => r := x"3ed3c2fd3fa4a331";
      when 1137 => r := x"3ed3a0f53fa495f6";
      when 1138 => r := x"3ed37ef63fa488bd";
      when 1139 => r := x"3ed35cfe3fa47b86";
      when 1140 => r := x"3ed33b0f3fa46e51";
      when 1141 => r := x"3ed319283fa4611f";
      when 1142 => r := x"3ed2f7493fa453ee";
      when 1143 => r := x"3ed2d5723fa446c0";
      when 1144 => r := x"3ed2b3a33fa43993";
      when 1145 => r := x"3ed291dd3fa42c69";
      when 1146 => r := x"3ed2701e3fa41f41";
      when 1147 => r := x"3ed24e683fa4121b";
      when 1148 => r := x"3ed22cba3fa404f7";
      when 1149 => r := x"3ed20b143fa3f7d6";
      when 1150 => r := x"3ed1e9763fa3eab6";
      when 1151 => r := x"3ed1c7e03fa3dd98";
      when 1152 => r := x"3ed1a6523fa3d07d";
      when 1153 => r := x"3ed184cc3fa3c364";
      when 1154 => r := x"3ed1634e3fa3b64c";
      when 1155 => r := x"3ed141d83fa3a937";
      when 1156 => r := x"3ed1206a3fa39c24";
      when 1157 => r := x"3ed0ff053fa38f13";
      when 1158 => r := x"3ed0dda73fa38204";
      when 1159 => r := x"3ed0bc513fa374f7";
      when 1160 => r := x"3ed09b033fa367ed";
      when 1161 => r := x"3ed079bd3fa35ae4";
      when 1162 => r := x"3ed0587f3fa34dde";
      when 1163 => r := x"3ed037493fa340d9";
      when 1164 => r := x"3ed0161b3fa333d7";
      when 1165 => r := x"3ecff4f53fa326d6";
      when 1166 => r := x"3ecfd3d73fa319d8";
      when 1167 => r := x"3ecfb2c13fa30cdc";
      when 1168 => r := x"3ecf91b23fa2ffe2";
      when 1169 => r := x"3ecf70ac3fa2f2ea";
      when 1170 => r := x"3ecf4fad3fa2e5f4";
      when 1171 => r := x"3ecf2eb73fa2d900";
      when 1172 => r := x"3ecf0dc83fa2cc0e";
      when 1173 => r := x"3eceece13fa2bf1e";
      when 1174 => r := x"3ececc023fa2b230";
      when 1175 => r := x"3eceab2a3fa2a544";
      when 1176 => r := x"3ece8a5b3fa2985b";
      when 1177 => r := x"3ece69933fa28b73";
      when 1178 => r := x"3ece48d33fa27e8e";
      when 1179 => r := x"3ece281b3fa271aa";
      when 1180 => r := x"3ece076b3fa264c8";
      when 1181 => r := x"3ecde6c23fa257e9";
      when 1182 => r := x"3ecdc6213fa24b0c";
      when 1183 => r := x"3ecda5883fa23e30";
      when 1184 => r := x"3ecd84f73fa23157";
      when 1185 => r := x"3ecd646d3fa22480";
      when 1186 => r := x"3ecd43ec3fa217aa";
      when 1187 => r := x"3ecd23713fa20ad7";
      when 1188 => r := x"3ecd02ff3fa1fe06";
      when 1189 => r := x"3ecce2943fa1f137";
      when 1190 => r := x"3eccc2313fa1e46a";
      when 1191 => r := x"3ecca1d63fa1d79f";
      when 1192 => r := x"3ecc81823fa1cad5";
      when 1193 => r := x"3ecc61363fa1be0e";
      when 1194 => r := x"3ecc40f23fa1b149";
      when 1195 => r := x"3ecc20b53fa1a486";
      when 1196 => r := x"3ecc00803fa197c5";
      when 1197 => r := x"3ecbe0523fa18b06";
      when 1198 => r := x"3ecbc02c3fa17e49";
      when 1199 => r := x"3ecba00e3fa1718e";
      when 1200 => r := x"3ecb7ff73fa164d5";
      when 1201 => r := x"3ecb5fe83fa1581e";
      when 1202 => r := x"3ecb3fe13fa14b69";
      when 1203 => r := x"3ecb1fe13fa13eb6";
      when 1204 => r := x"3ecaffe83fa13205";
      when 1205 => r := x"3ecadff73fa12556";
      when 1206 => r := x"3ecac00e3fa118a9";
      when 1207 => r := x"3ecaa02c3fa10bfe";
      when 1208 => r := x"3eca80523fa0ff55";
      when 1209 => r := x"3eca607f3fa0f2ae";
      when 1210 => r := x"3eca40b43fa0e609";
      when 1211 => r := x"3eca20f03fa0d966";
      when 1212 => r := x"3eca01343fa0ccc5";
      when 1213 => r := x"3ec9e17f3fa0c026";
      when 1214 => r := x"3ec9c1d23fa0b389";
      when 1215 => r := x"3ec9a22c3fa0a6ee";
      when 1216 => r := x"3ec9828d3fa09a54";
      when 1217 => r := x"3ec962f63fa08dbd";
      when 1218 => r := x"3ec943663fa08128";
      when 1219 => r := x"3ec923de3fa07495";
      when 1220 => r := x"3ec9045d3fa06804";
      when 1221 => r := x"3ec8e4e43fa05b74";
      when 1222 => r := x"3ec8c5723fa04ee7";
      when 1223 => r := x"3ec8a6073fa0425c";
      when 1224 => r := x"3ec886a43fa035d2";
      when 1225 => r := x"3ec867483fa0294b";
      when 1226 => r := x"3ec847f43fa01cc5";
      when 1227 => r := x"3ec828a63fa01042";
      when 1228 => r := x"3ec809613fa003c0";
      when 1229 => r := x"3ec7ea223f9ff741";
      when 1230 => r := x"3ec7caeb3f9feac3";
      when 1231 => r := x"3ec7abbb3f9fde47";
      when 1232 => r := x"3ec78c923f9fd1ce";
      when 1233 => r := x"3ec76d713f9fc556";
      when 1234 => r := x"3ec74e573f9fb8e0";
      when 1235 => r := x"3ec72f443f9fac6c";
      when 1236 => r := x"3ec710393f9f9ffa";
      when 1237 => r := x"3ec6f1353f9f938a";
      when 1238 => r := x"3ec6d2383f9f871c";
      when 1239 => r := x"3ec6b3423f9f7ab0";
      when 1240 => r := x"3ec694533f9f6e45";
      when 1241 => r := x"3ec6756c3f9f61dd";
      when 1242 => r := x"3ec6568c3f9f5577";
      when 1243 => r := x"3ec637b33f9f4912";
      when 1244 => r := x"3ec618e13f9f3cb0";
      when 1245 => r := x"3ec5fa173f9f304f";
      when 1246 => r := x"3ec5db533f9f23f0";
      when 1247 => r := x"3ec5bc973f9f1794";
      when 1248 => r := x"3ec59de23f9f0b39";
      when 1249 => r := x"3ec57f343f9efee0";
      when 1250 => r := x"3ec5608e3f9ef289";
      when 1251 => r := x"3ec541ee3f9ee634";
      when 1252 => r := x"3ec523563f9ed9e1";
      when 1253 => r := x"3ec504c43f9ecd90";
      when 1254 => r := x"3ec4e63a3f9ec140";
      when 1255 => r := x"3ec4c7b73f9eb4f3";
      when 1256 => r := x"3ec4a93b3f9ea8a7";
      when 1257 => r := x"3ec48ac63f9e9c5e";
      when 1258 => r := x"3ec46c583f9e9016";
      when 1259 => r := x"3ec44df13f9e83d0";
      when 1260 => r := x"3ec42f913f9e778c";
      when 1261 => r := x"3ec411393f9e6b4a";
      when 1262 => r := x"3ec3f2e73f9e5f0a";
      when 1263 => r := x"3ec3d49c3f9e52cc";
      when 1264 => r := x"3ec3b6593f9e468f";
      when 1265 => r := x"3ec3981c3f9e3a55";
      when 1266 => r := x"3ec379e63f9e2e1c";
      when 1267 => r := x"3ec35bb83f9e21e6";
      when 1268 => r := x"3ec33d903f9e15b1";
      when 1269 => r := x"3ec31f703f9e097e";
      when 1270 => r := x"3ec301563f9dfd4d";
      when 1271 => r := x"3ec2e3433f9df11e";
      when 1272 => r := x"3ec2c5373f9de4f1";
      when 1273 => r := x"3ec2a7333f9dd8c5";
      when 1274 => r := x"3ec289353f9dcc9c";
      when 1275 => r := x"3ec26b3e3f9dc074";
      when 1276 => r := x"3ec24d4e3f9db44e";
      when 1277 => r := x"3ec22f653f9da82a";
      when 1278 => r := x"3ec211833f9d9c08";
      when 1279 => r := x"3ec1f3a73f9d8fe8";
      when 1280 => r := x"3ec1d5d33f9d83ca";
      when 1281 => r := x"3ec1b8053f9d77ad";
      when 1282 => r := x"3ec19a3f3f9d6b93";
      when 1283 => r := x"3ec17c7f3f9d5f7a";
      when 1284 => r := x"3ec15ec63f9d5363";
      when 1285 => r := x"3ec141143f9d474e";
      when 1286 => r := x"3ec123683f9d3b3b";
      when 1287 => r := x"3ec105c43f9d2f2a";
      when 1288 => r := x"3ec0e8263f9d231a";
      when 1289 => r := x"3ec0ca903f9d170d";
      when 1290 => r := x"3ec0ad003f9d0b01";
      when 1291 => r := x"3ec08f763f9cfef7";
      when 1292 => r := x"3ec071f43f9cf2ef";
      when 1293 => r := x"3ec054783f9ce6e9";
      when 1294 => r := x"3ec037033f9cdae5";
      when 1295 => r := x"3ec019953f9ccee2";
      when 1296 => r := x"3ebffc2e3f9cc2e1";
      when 1297 => r := x"3ebfdecd3f9cb6e3";
      when 1298 => r := x"3ebfc1743f9caae6";
      when 1299 => r := x"3ebfa4213f9c9eea";
      when 1300 => r := x"3ebf86d43f9c92f1";
      when 1301 => r := x"3ebf698e3f9c86fa";
      when 1302 => r := x"3ebf4c503f9c7b04";
      when 1303 => r := x"3ebf2f173f9c6f10";
      when 1304 => r := x"3ebf11e63f9c631e";
      when 1305 => r := x"3ebef4bb3f9c572e";
      when 1306 => r := x"3ebed7973f9c4b3f";
      when 1307 => r := x"3ebeba793f9c3f53";
      when 1308 => r := x"3ebe9d623f9c3368";
      when 1309 => r := x"3ebe80523f9c277f";
      when 1310 => r := x"3ebe63483f9c1b98";
      when 1311 => r := x"3ebe46453f9c0fb3";
      when 1312 => r := x"3ebe29493f9c03cf";
      when 1313 => r := x"3ebe0c533f9bf7ee";
      when 1314 => r := x"3ebdef643f9bec0e";
      when 1315 => r := x"3ebdd27c3f9be030";
      when 1316 => r := x"3ebdb59a3f9bd453";
      when 1317 => r := x"3ebd98bf3f9bc879";
      when 1318 => r := x"3ebd7bea3f9bbca0";
      when 1319 => r := x"3ebd5f1c3f9bb0c9";
      when 1320 => r := x"3ebd42543f9ba4f4";
      when 1321 => r := x"3ebd25933f9b9921";
      when 1322 => r := x"3ebd08d93f9b8d50";
      when 1323 => r := x"3ebcec253f9b8180";
      when 1324 => r := x"3ebccf783f9b75b2";
      when 1325 => r := x"3ebcb2d13f9b69e6";
      when 1326 => r := x"3ebc96313f9b5e1c";
      when 1327 => r := x"3ebc79973f9b5253";
      when 1328 => r := x"3ebc5d033f9b468d";
      when 1329 => r := x"3ebc40773f9b3ac8";
      when 1330 => r := x"3ebc23f03f9b2f05";
      when 1331 => r := x"3ebc07703f9b2343";
      when 1332 => r := x"3ebbeaf73f9b1784";
      when 1333 => r := x"3ebbce843f9b0bc6";
      when 1334 => r := x"3ebbb2183f9b000a";
      when 1335 => r := x"3ebb95b23f9af450";
      when 1336 => r := x"3ebb79523f9ae897";
      when 1337 => r := x"3ebb5cf93f9adce0";
      when 1338 => r := x"3ebb40a63f9ad12c";
      when 1339 => r := x"3ebb245a3f9ac578";
      when 1340 => r := x"3ebb08143f9ab9c7";
      when 1341 => r := x"3ebaebd53f9aae17";
      when 1342 => r := x"3ebacf9c3f9aa269";
      when 1343 => r := x"3ebab3693f9a96bd";
      when 1344 => r := x"3eba973d3f9a8b13";
      when 1345 => r := x"3eba7b173f9a7f6a";
      when 1346 => r := x"3eba5ef73f9a73c4";
      when 1347 => r := x"3eba42de3f9a681f";
      when 1348 => r := x"3eba26cb3f9a5c7b";
      when 1349 => r := x"3eba0abf3f9a50da";
      when 1350 => r := x"3eb9eeb93f9a453a";
      when 1351 => r := x"3eb9d2b93f9a399c";
      when 1352 => r := x"3eb9b6c03f9a2e00";
      when 1353 => r := x"3eb99acc3f9a2265";
      when 1354 => r := x"3eb97edf3f9a16cc";
      when 1355 => r := x"3eb962f93f9a0b35";
      when 1356 => r := x"3eb947193f99ffa0";
      when 1357 => r := x"3eb92b3f3f99f40c";
      when 1358 => r := x"3eb90f6b3f99e87b";
      when 1359 => r := x"3eb8f39e3f99dcea";
      when 1360 => r := x"3eb8d7d63f99d15c";
      when 1361 => r := x"3eb8bc153f99c5cf";
      when 1362 => r := x"3eb8a05b3f99ba45";
      when 1363 => r := x"3eb884a63f99aebb";
      when 1364 => r := x"3eb868f83f99a334";
      when 1365 => r := x"3eb84d503f9997ae";
      when 1366 => r := x"3eb831ae3f998c2a";
      when 1367 => r := x"3eb816133f9980a8";
      when 1368 => r := x"3eb7fa7e3f997528";
      when 1369 => r := x"3eb7deee3f9969a9";
      when 1370 => r := x"3eb7c3663f995e2c";
      when 1371 => r := x"3eb7a7e33f9952b0";
      when 1372 => r := x"3eb78c663f994737";
      when 1373 => r := x"3eb770f03f993bbf";
      when 1374 => r := x"3eb755803f993049";
      when 1375 => r := x"3eb73a153f9924d4";
      when 1376 => r := x"3eb71eb23f991961";
      when 1377 => r := x"3eb703543f990df0";
      when 1378 => r := x"3eb6e7fc3f990281";
      when 1379 => r := x"3eb6ccaa3f98f713";
      when 1380 => r := x"3eb6b15f3f98eba7";
      when 1381 => r := x"3eb6961a3f98e03d";
      when 1382 => r := x"3eb67adb3f98d4d5";
      when 1383 => r := x"3eb65fa13f98c96e";
      when 1384 => r := x"3eb6446e3f98be09";
      when 1385 => r := x"3eb629413f98b2a5";
      when 1386 => r := x"3eb60e1b3f98a743";
      when 1387 => r := x"3eb5f2fa3f989be3";
      when 1388 => r := x"3eb5d7df3f989085";
      when 1389 => r := x"3eb5bcca3f988528";
      when 1390 => r := x"3eb5a1bc3f9879cd";
      when 1391 => r := x"3eb586b33f986e74";
      when 1392 => r := x"3eb56bb13f98631d";
      when 1393 => r := x"3eb550b43f9857c7";
      when 1394 => r := x"3eb535be3f984c73";
      when 1395 => r := x"3eb51acd3f984120";
      when 1396 => r := x"3eb4ffe33f9835cf";
      when 1397 => r := x"3eb4e4fe3f982a80";
      when 1398 => r := x"3eb4ca203f981f33";
      when 1399 => r := x"3eb4af473f9813e7";
      when 1400 => r := x"3eb494743f98089d";
      when 1401 => r := x"3eb479a83f97fd54";
      when 1402 => r := x"3eb45ee13f97f20d";
      when 1403 => r := x"3eb444213f97e6c8";
      when 1404 => r := x"3eb429663f97db85";
      when 1405 => r := x"3eb40eb13f97d043";
      when 1406 => r := x"3eb3f4023f97c503";
      when 1407 => r := x"3eb3d9593f97b9c5";
      when 1408 => r := x"3eb3beb73f97ae88";
      when 1409 => r := x"3eb3a4193f97a34d";
      when 1410 => r := x"3eb389823f979813";
      when 1411 => r := x"3eb36ef13f978cdc";
      when 1412 => r := x"3eb354663f9781a6";
      when 1413 => r := x"3eb339e03f977671";
      when 1414 => r := x"3eb31f613f976b3e";
      when 1415 => r := x"3eb304e73f97600d";
      when 1416 => r := x"3eb2ea733f9754de";
      when 1417 => r := x"3eb2d0053f9749b0";
      when 1418 => r := x"3eb2b59d3f973e84";
      when 1419 => r := x"3eb29b3b3f973359";
      when 1420 => r := x"3eb280de3f972830";
      when 1421 => r := x"3eb266883f971d09";
      when 1422 => r := x"3eb24c373f9711e3";
      when 1423 => r := x"3eb231ec3f9706c0";
      when 1424 => r := x"3eb217a73f96fb9d";
      when 1425 => r := x"3eb1fd683f96f07d";
      when 1426 => r := x"3eb1e32e3f96e55e";
      when 1427 => r := x"3eb1c8fa3f96da40";
      when 1428 => r := x"3eb1aecc3f96cf24";
      when 1429 => r := x"3eb194a43f96c40a";
      when 1430 => r := x"3eb17a823f96b8f2";
      when 1431 => r := x"3eb160653f96addb";
      when 1432 => r := x"3eb1464e3f96a2c6";
      when 1433 => r := x"3eb12c3d3f9697b2";
      when 1434 => r := x"3eb112323f968ca0";
      when 1435 => r := x"3eb0f82c3f968190";
      when 1436 => r := x"3eb0de2c3f967681";
      when 1437 => r := x"3eb0c4323f966b74";
      when 1438 => r := x"3eb0aa3e3f966069";
      when 1439 => r := x"3eb0904f3f96555f";
      when 1440 => r := x"3eb076663f964a57";
      when 1441 => r := x"3eb05c833f963f50";
      when 1442 => r := x"3eb042a53f96344b";
      when 1443 => r := x"3eb028cd3f962948";
      when 1444 => r := x"3eb00efb3f961e46";
      when 1445 => r := x"3eaff52f3f961346";
      when 1446 => r := x"3eafdb683f960847";
      when 1447 => r := x"3eafc1a63f95fd4a";
      when 1448 => r := x"3eafa7eb3f95f24f";
      when 1449 => r := x"3eaf8e353f95e755";
      when 1450 => r := x"3eaf74853f95dc5d";
      when 1451 => r := x"3eaf5ada3f95d167";
      when 1452 => r := x"3eaf41353f95c672";
      when 1453 => r := x"3eaf27963f95bb7f";
      when 1454 => r := x"3eaf0dfc3f95b08d";
      when 1455 => r := x"3eaef4683f95a59d";
      when 1456 => r := x"3eaedad93f959aaf";
      when 1457 => r := x"3eaec1503f958fc2";
      when 1458 => r := x"3eaea7cd3f9584d6";
      when 1459 => r := x"3eae8e4f3f9579ed";
      when 1460 => r := x"3eae74d73f956f05";
      when 1461 => r := x"3eae5b643f95641e";
      when 1462 => r := x"3eae41f73f955939";
      when 1463 => r := x"3eae28903f954e56";
      when 1464 => r := x"3eae0f2e3f954374";
      when 1465 => r := x"3eadf5d13f953894";
      when 1466 => r := x"3eaddc7a3f952db5";
      when 1467 => r := x"3eadc3293f9522d8";
      when 1468 => r := x"3eada9dd3f9517fd";
      when 1469 => r := x"3ead90973f950d23";
      when 1470 => r := x"3ead77563f95024b";
      when 1471 => r := x"3ead5e1b3f94f774";
      when 1472 => r := x"3ead44e53f94ec9f";
      when 1473 => r := x"3ead2bb53f94e1cc";
      when 1474 => r := x"3ead128a3f94d6fa";
      when 1475 => r := x"3eacf9653f94cc29";
      when 1476 => r := x"3eace0453f94c15a";
      when 1477 => r := x"3eacc72b3f94b68d";
      when 1478 => r := x"3eacae163f94abc2";
      when 1479 => r := x"3eac95073f94a0f7";
      when 1480 => r := x"3eac7bfd3f94962f";
      when 1481 => r := x"3eac62f83f948b68";
      when 1482 => r := x"3eac49f93f9480a3";
      when 1483 => r := x"3eac30ff3f9475df";
      when 1484 => r := x"3eac180b3f946b1c";
      when 1485 => r := x"3eabff1d3f94605c";
      when 1486 => r := x"3eabe6333f94559d";
      when 1487 => r := x"3eabcd4f3f944adf";
      when 1488 => r := x"3eabb4713f944023";
      when 1489 => r := x"3eab9b983f943568";
      when 1490 => r := x"3eab82c43f942aaf";
      when 1491 => r := x"3eab69f53f941ff8";
      when 1492 => r := x"3eab512c3f941542";
      when 1493 => r := x"3eab38693f940a8e";
      when 1494 => r := x"3eab1fab3f93ffdb";
      when 1495 => r := x"3eab06f23f93f52a";
      when 1496 => r := x"3eaaee3e3f93ea7a";
      when 1497 => r := x"3eaad5903f93dfcc";
      when 1498 => r := x"3eaabce73f93d520";
      when 1499 => r := x"3eaaa4443f93ca75";
      when 1500 => r := x"3eaa8ba63f93bfcb";
      when 1501 => r := x"3eaa730d3f93b523";
      when 1502 => r := x"3eaa5a793f93aa7d";
      when 1503 => r := x"3eaa41eb3f939fd8";
      when 1504 => r := x"3eaa29623f939534";
      when 1505 => r := x"3eaa10df3f938a93";
      when 1506 => r := x"3ea9f8603f937ff2";
      when 1507 => r := x"3ea9dfe73f937554";
      when 1508 => r := x"3ea9c7743f936ab6";
      when 1509 => r := x"3ea9af053f93601b";
      when 1510 => r := x"3ea9969c3f935580";
      when 1511 => r := x"3ea97e383f934ae8";
      when 1512 => r := x"3ea965d93f934051";
      when 1513 => r := x"3ea94d803f9335bb";
      when 1514 => r := x"3ea9352c3f932b27";
      when 1515 => r := x"3ea91cdd3f932094";
      when 1516 => r := x"3ea904933f931603";
      when 1517 => r := x"3ea8ec4f3f930b74";
      when 1518 => r := x"3ea8d4103f9300e6";
      when 1519 => r := x"3ea8bbd63f92f659";
      when 1520 => r := x"3ea8a3a13f92ebce";
      when 1521 => r := x"3ea88b713f92e145";
      when 1522 => r := x"3ea873473f92d6bd";
      when 1523 => r := x"3ea85b223f92cc36";
      when 1524 => r := x"3ea843023f92c1b2";
      when 1525 => r := x"3ea82ae73f92b72e";
      when 1526 => r := x"3ea812d23f92acac";
      when 1527 => r := x"3ea7fac13f92a22c";
      when 1528 => r := x"3ea7e2b63f9297ad";
      when 1529 => r := x"3ea7cab03f928d2f";
      when 1530 => r := x"3ea7b2af3f9282b3";
      when 1531 => r := x"3ea79ab33f927839";
      when 1532 => r := x"3ea782bc3f926dc0";
      when 1533 => r := x"3ea76acb3f926349";
      when 1534 => r := x"3ea752de3f9258d3";
      when 1535 => r := x"3ea73af73f924e5e";
      when 1536 => r := x"3ea723153f9243eb";
      when 1537 => r := x"3ea70b383f92397a";
      when 1538 => r := x"3ea6f3603f922f0a";
      when 1539 => r := x"3ea6db8d3f92249c";
      when 1540 => r := x"3ea6c3c03f921a2f";
      when 1541 => r := x"3ea6abf73f920fc3";
      when 1542 => r := x"3ea694333f920559";
      when 1543 => r := x"3ea67c753f91faf1";
      when 1544 => r := x"3ea664bb3f91f08a";
      when 1545 => r := x"3ea64d073f91e624";
      when 1546 => r := x"3ea635583f91dbc0";
      when 1547 => r := x"3ea61dae3f91d15d";
      when 1548 => r := x"3ea606093f91c6fc";
      when 1549 => r := x"3ea5ee693f91bc9d";
      when 1550 => r := x"3ea5d6cd3f91b23e";
      when 1551 => r := x"3ea5bf373f91a7e2";
      when 1552 => r := x"3ea5a7a63f919d86";
      when 1553 => r := x"3ea5901a3f91932d";
      when 1554 => r := x"3ea578943f9188d4";
      when 1555 => r := x"3ea561123f917e7e";
      when 1556 => r := x"3ea549953f917428";
      when 1557 => r := x"3ea5321d3f9169d4";
      when 1558 => r := x"3ea51aaa3f915f82";
      when 1559 => r := x"3ea5033c3f915531";
      when 1560 => r := x"3ea4ebd33f914ae2";
      when 1561 => r := x"3ea4d46f3f914094";
      when 1562 => r := x"3ea4bd103f913647";
      when 1563 => r := x"3ea4a5b63f912bfc";
      when 1564 => r := x"3ea48e613f9121b2";
      when 1565 => r := x"3ea477113f91176a";
      when 1566 => r := x"3ea45fc63f910d24";
      when 1567 => r := x"3ea448803f9102de";
      when 1568 => r := x"3ea4313e3f90f89a";
      when 1569 => r := x"3ea41a023f90ee58";
      when 1570 => r := x"3ea402cb3f90e417";
      when 1571 => r := x"3ea3eb983f90d9d8";
      when 1572 => r := x"3ea3d46b3f90cf9a";
      when 1573 => r := x"3ea3bd423f90c55d";
      when 1574 => r := x"3ea3a61e3f90bb22";
      when 1575 => r := x"3ea38eff3f90b0e8";
      when 1576 => r := x"3ea377e53f90a6b0";
      when 1577 => r := x"3ea360d03f909c79";
      when 1578 => r := x"3ea349c03f909244";
      when 1579 => r := x"3ea332b53f908810";
      when 1580 => r := x"3ea31baf3f907dde";
      when 1581 => r := x"3ea304ad3f9073ad";
      when 1582 => r := x"3ea2edb13f90697d";
      when 1583 => r := x"3ea2d6b93f905f4f";
      when 1584 => r := x"3ea2bfc63f905522";
      when 1585 => r := x"3ea2a8d83f904af7";
      when 1586 => r := x"3ea291ef3f9040cd";
      when 1587 => r := x"3ea27b0a3f9036a5";
      when 1588 => r := x"3ea2642b3f902c7e";
      when 1589 => r := x"3ea24d503f902258";
      when 1590 => r := x"3ea2367a3f901834";
      when 1591 => r := x"3ea21fa93f900e12";
      when 1592 => r := x"3ea208dd3f9003f0";
      when 1593 => r := x"3ea1f2153f8ff9d0";
      when 1594 => r := x"3ea1db523f8fefb2";
      when 1595 => r := x"3ea1c4953f8fe595";
      when 1596 => r := x"3ea1addb3f8fdb79";
      when 1597 => r := x"3ea197273f8fd15f";
      when 1598 => r := x"3ea180783f8fc747";
      when 1599 => r := x"3ea169cd3f8fbd2f";
      when 1600 => r := x"3ea153273f8fb319";
      when 1601 => r := x"3ea13c863f8fa905";
      when 1602 => r := x"3ea125e93f8f9ef2";
      when 1603 => r := x"3ea10f523f8f94e0";
      when 1604 => r := x"3ea0f8bf3f8f8ad0";
      when 1605 => r := x"3ea0e2313f8f80c1";
      when 1606 => r := x"3ea0cba73f8f76b4";
      when 1607 => r := x"3ea0b5223f8f6ca8";
      when 1608 => r := x"3ea09ea23f8f629d";
      when 1609 => r := x"3ea088273f8f5894";
      when 1610 => r := x"3ea071b13f8f4e8c";
      when 1611 => r := x"3ea05b3f3f8f4485";
      when 1612 => r := x"3ea044d23f8f3a80";
      when 1613 => r := x"3ea02e693f8f307d";
      when 1614 => r := x"3ea018063f8f267b";
      when 1615 => r := x"3ea001a73f8f1c7a";
      when 1616 => r := x"3e9feb4c3f8f127a";
      when 1617 => r := x"3e9fd4f73f8f087c";
      when 1618 => r := x"3e9fbea63f8efe80";
      when 1619 => r := x"3e9fa8593f8ef485";
      when 1620 => r := x"3e9f92123f8eea8b";
      when 1621 => r := x"3e9f7bcf3f8ee092";
      when 1622 => r := x"3e9f65903f8ed69b";
      when 1623 => r := x"3e9f4f573f8ecca6";
      when 1624 => r := x"3e9f39223f8ec2b1";
      when 1625 => r := x"3e9f22f13f8eb8bf";
      when 1626 => r := x"3e9f0cc63f8eaecd";
      when 1627 => r := x"3e9ef69e3f8ea4dd";
      when 1628 => r := x"3e9ee07c3f8e9aee";
      when 1629 => r := x"3e9eca5e3f8e9101";
      when 1630 => r := x"3e9eb4453f8e8715";
      when 1631 => r := x"3e9e9e303f8e7d2a";
      when 1632 => r := x"3e9e88203f8e7341";
      when 1633 => r := x"3e9e72153f8e6959";
      when 1634 => r := x"3e9e5c0e3f8e5f73";
      when 1635 => r := x"3e9e460c3f8e558e";
      when 1636 => r := x"3e9e300e3f8e4baa";
      when 1637 => r := x"3e9e1a153f8e41c8";
      when 1638 => r := x"3e9e04213f8e37e7";
      when 1639 => r := x"3e9dee313f8e2e07";
      when 1640 => r := x"3e9dd8453f8e2429";
      when 1641 => r := x"3e9dc25e3f8e1a4c";
      when 1642 => r := x"3e9dac7c3f8e1071";
      when 1643 => r := x"3e9d969f3f8e0697";
      when 1644 => r := x"3e9d80c53f8dfcbe";
      when 1645 => r := x"3e9d6af13f8df2e7";
      when 1646 => r := x"3e9d55213f8de911";
      when 1647 => r := x"3e9d3f553f8ddf3c";
      when 1648 => r := x"3e9d298e3f8dd569";
      when 1649 => r := x"3e9d13cc3f8dcb97";
      when 1650 => r := x"3e9cfe0e3f8dc1c6";
      when 1651 => r := x"3e9ce8543f8db7f7";
      when 1652 => r := x"3e9cd2a03f8dae29";
      when 1653 => r := x"3e9cbcef3f8da45d";
      when 1654 => r := x"3e9ca7433f8d9a92";
      when 1655 => r := x"3e9c919c3f8d90c8";
      when 1656 => r := x"3e9c7bf93f8d86ff";
      when 1657 => r := x"3e9c665a3f8d7d38";
      when 1658 => r := x"3e9c50c03f8d7373";
      when 1659 => r := x"3e9c3b2b3f8d69ae";
      when 1660 => r := x"3e9c259a3f8d5feb";
      when 1661 => r := x"3e9c100d3f8d5629";
      when 1662 => r := x"3e9bfa853f8d4c69";
      when 1663 => r := x"3e9be5013f8d42aa";
      when 1664 => r := x"3e9bcf823f8d38ed";
      when 1665 => r := x"3e9bba083f8d2f30";
      when 1666 => r := x"3e9ba4913f8d2575";
      when 1667 => r := x"3e9b8f1f3f8d1bbc";
      when 1668 => r := x"3e9b79b23f8d1203";
      when 1669 => r := x"3e9b64493f8d084c";
      when 1670 => r := x"3e9b4ee43f8cfe97";
      when 1671 => r := x"3e9b39843f8cf4e3";
      when 1672 => r := x"3e9b24283f8ceb30";
      when 1673 => r := x"3e9b0ed13f8ce17e";
      when 1674 => r := x"3e9af97e3f8cd7ce";
      when 1675 => r := x"3e9ae42f3f8cce1f";
      when 1676 => r := x"3e9acee53f8cc471";
      when 1677 => r := x"3e9ab99f3f8cbac5";
      when 1678 => r := x"3e9aa45e3f8cb11a";
      when 1679 => r := x"3e9a8f213f8ca770";
      when 1680 => r := x"3e9a79e83f8c9dc8";
      when 1681 => r := x"3e9a64b43f8c9421";
      when 1682 => r := x"3e9a4f843f8c8a7c";
      when 1683 => r := x"3e9a3a583f8c80d7";
      when 1684 => r := x"3e9a25313f8c7734";
      when 1685 => r := x"3e9a100e3f8c6d93";
      when 1686 => r := x"3e99faf03f8c63f2";
      when 1687 => r := x"3e99e5d63f8c5a53";
      when 1688 => r := x"3e99d0c03f8c50b6";
      when 1689 => r := x"3e99bbae3f8c4719";
      when 1690 => r := x"3e99a6a13f8c3d7e";
      when 1691 => r := x"3e9991983f8c33e4";
      when 1692 => r := x"3e997c943f8c2a4c";
      when 1693 => r := x"3e9967943f8c20b5";
      when 1694 => r := x"3e9952983f8c171f";
      when 1695 => r := x"3e993da03f8c0d8a";
      when 1696 => r := x"3e9928ad3f8c03f7";
      when 1697 => r := x"3e9913be3f8bfa65";
      when 1698 => r := x"3e98fed33f8bf0d5";
      when 1699 => r := x"3e98e9ed3f8be745";
      when 1700 => r := x"3e98d50b3f8bddb8";
      when 1701 => r := x"3e98c02d3f8bd42b";
      when 1702 => r := x"3e98ab533f8bcaa0";
      when 1703 => r := x"3e98967e3f8bc115";
      when 1704 => r := x"3e9881ad3f8bb78d";
      when 1705 => r := x"3e986ce03f8bae05";
      when 1706 => r := x"3e9858173f8ba47f";
      when 1707 => r := x"3e9843533f8b9afa";
      when 1708 => r := x"3e982e933f8b9177";
      when 1709 => r := x"3e9819d73f8b87f4";
      when 1710 => r := x"3e9805203f8b7e73";
      when 1711 => r := x"3e97f06c3f8b74f4";
      when 1712 => r := x"3e97dbbd3f8b6b75";
      when 1713 => r := x"3e97c7123f8b61f8";
      when 1714 => r := x"3e97b26b3f8b587c";
      when 1715 => r := x"3e979dc93f8b4f02";
      when 1716 => r := x"3e97892b3f8b4589";
      when 1717 => r := x"3e9774913f8b3c11";
      when 1718 => r := x"3e975ffb3f8b329a";
      when 1719 => r := x"3e974b693f8b2925";
      when 1720 => r := x"3e9736dc3f8b1fb1";
      when 1721 => r := x"3e9722523f8b163e";
      when 1722 => r := x"3e970dcd3f8b0ccc";
      when 1723 => r := x"3e96f94c3f8b035c";
      when 1724 => r := x"3e96e4d03f8af9ed";
      when 1725 => r := x"3e96d0573f8af080";
      when 1726 => r := x"3e96bbe33f8ae713";
      when 1727 => r := x"3e96a7723f8adda8";
      when 1728 => r := x"3e9693063f8ad43e";
      when 1729 => r := x"3e967e9e3f8acad6";
      when 1730 => r := x"3e966a3b3f8ac16f";
      when 1731 => r := x"3e9655db3f8ab809";
      when 1732 => r := x"3e96417f3f8aaea4";
      when 1733 => r := x"3e962d283f8aa540";
      when 1734 => r := x"3e9618d53f8a9bde";
      when 1735 => r := x"3e9604863f8a927d";
      when 1736 => r := x"3e95f03b3f8a891e";
      when 1737 => r := x"3e95dbf43f8a7fbf";
      when 1738 => r := x"3e95c7b13f8a7662";
      when 1739 => r := x"3e95b3723f8a6d06";
      when 1740 => r := x"3e959f383f8a63ac";
      when 1741 => r := x"3e958b013f8a5a52";
      when 1742 => r := x"3e9576cf3f8a50fa";
      when 1743 => r := x"3e9562a13f8a47a3";
      when 1744 => r := x"3e954e763f8a3e4e";
      when 1745 => r := x"3e953a503f8a34fa";
      when 1746 => r := x"3e95262e3f8a2ba7";
      when 1747 => r := x"3e9512103f8a2255";
      when 1748 => r := x"3e94fdf63f8a1904";
      when 1749 => r := x"3e94e9e03f8a0fb5";
      when 1750 => r := x"3e94d5cf3f8a0667";
      when 1751 => r := x"3e94c1c13f89fd1a";
      when 1752 => r := x"3e94adb73f89f3cf";
      when 1753 => r := x"3e9499b23f89ea85";
      when 1754 => r := x"3e9485b03f89e13c";
      when 1755 => r := x"3e9471b33f89d7f4";
      when 1756 => r := x"3e945db93f89ceae";
      when 1757 => r := x"3e9449c43f89c568";
      when 1758 => r := x"3e9435d23f89bc24";
      when 1759 => r := x"3e9421e53f89b2e2";
      when 1760 => r := x"3e940dfb3f89a9a0";
      when 1761 => r := x"3e93fa163f89a060";
      when 1762 => r := x"3e93e6353f899721";
      when 1763 => r := x"3e93d2573f898de3";
      when 1764 => r := x"3e93be7e3f8984a7";
      when 1765 => r := x"3e93aaa83f897b6b";
      when 1766 => r := x"3e9396d73f897231";
      when 1767 => r := x"3e93830a3f8968f8";
      when 1768 => r := x"3e936f403f895fc1";
      when 1769 => r := x"3e935b7b3f89568a";
      when 1770 => r := x"3e9347b93f894d55";
      when 1771 => r := x"3e9333fc3f894421";
      when 1772 => r := x"3e9320423f893aef";
      when 1773 => r := x"3e930c8d3f8931bd";
      when 1774 => r := x"3e92f8db3f89288d";
      when 1775 => r := x"3e92e52e3f891f5e";
      when 1776 => r := x"3e92d1843f891631";
      when 1777 => r := x"3e92bdde3f890d04";
      when 1778 => r := x"3e92aa3c3f8903d9";
      when 1779 => r := x"3e92969e3f88faaf";
      when 1780 => r := x"3e9283053f88f186";
      when 1781 => r := x"3e926f6f3f88e85f";
      when 1782 => r := x"3e925bdd3f88df38";
      when 1783 => r := x"3e92484e3f88d613";
      when 1784 => r := x"3e9234c43f88ccef";
      when 1785 => r := x"3e92213e3f88c3cc";
      when 1786 => r := x"3e920dbb3f88baab";
      when 1787 => r := x"3e91fa3d3f88b18b";
      when 1788 => r := x"3e91e6c23f88a86c";
      when 1789 => r := x"3e91d34c3f889f4e";
      when 1790 => r := x"3e91bfd93f889631";
      when 1791 => r := x"3e91ac6a3f888d16";
      when 1792 => r := x"3e9198ff3f8883fc";
      when 1793 => r := x"3e9185983f887ae3";
      when 1794 => r := x"3e9172343f8871cb";
      when 1795 => r := x"3e915ed53f8868b4";
      when 1796 => r := x"3e914b7a3f885f9f";
      when 1797 => r := x"3e9138223f88568b";
      when 1798 => r := x"3e9124ce3f884d78";
      when 1799 => r := x"3e91117e3f884466";
      when 1800 => r := x"3e90fe323f883b56";
      when 1801 => r := x"3e90eaea3f883247";
      when 1802 => r := x"3e90d7a53f882939";
      when 1803 => r := x"3e90c4653f88202c";
      when 1804 => r := x"3e90b1283f881720";
      when 1805 => r := x"3e909def3f880e16";
      when 1806 => r := x"3e908aba3f88050c";
      when 1807 => r := x"3e9077893f87fc04";
      when 1808 => r := x"3e90645c3f87f2fd";
      when 1809 => r := x"3e9051323f87e9f8";
      when 1810 => r := x"3e903e0c3f87e0f3";
      when 1811 => r := x"3e902aea3f87d7f0";
      when 1812 => r := x"3e9017cc3f87ceee";
      when 1813 => r := x"3e9004b23f87c5ed";
      when 1814 => r := x"3e8ff19b3f87bced";
      when 1815 => r := x"3e8fde883f87b3ef";
      when 1816 => r := x"3e8fcb793f87aaf1";
      when 1817 => r := x"3e8fb86e3f87a1f5";
      when 1818 => r := x"3e8fa5673f8798fa";
      when 1819 => r := x"3e8f92633f879001";
      when 1820 => r := x"3e8f7f633f878708";
      when 1821 => r := x"3e8f6c673f877e11";
      when 1822 => r := x"3e8f596f3f87751b";
      when 1823 => r := x"3e8f467a3f876c26";
      when 1824 => r := x"3e8f338a3f876332";
      when 1825 => r := x"3e8f209d3f875a3f";
      when 1826 => r := x"3e8f0db33f87514e";
      when 1827 => r := x"3e8eface3f87485d";
      when 1828 => r := x"3e8ee7ec3f873f6e";
      when 1829 => r := x"3e8ed50e3f873680";
      when 1830 => r := x"3e8ec2343f872d94";
      when 1831 => r := x"3e8eaf5d3f8724a8";
      when 1832 => r := x"3e8e9c8a3f871bbe";
      when 1833 => r := x"3e8e89bb3f8712d5";
      when 1834 => r := x"3e8e76f03f8709ed";
      when 1835 => r := x"3e8e64283f870106";
      when 1836 => r := x"3e8e51643f86f820";
      when 1837 => r := x"3e8e3ea43f86ef3c";
      when 1838 => r := x"3e8e2be73f86e658";
      when 1839 => r := x"3e8e192e3f86dd76";
      when 1840 => r := x"3e8e06793f86d495";
      when 1841 => r := x"3e8df3c83f86cbb5";
      when 1842 => r := x"3e8de11a3f86c2d7";
      when 1843 => r := x"3e8dce703f86b9f9";
      when 1844 => r := x"3e8dbbc93f86b11d";
      when 1845 => r := x"3e8da9263f86a842";
      when 1846 => r := x"3e8d96873f869f68";
      when 1847 => r := x"3e8d83ec3f86968f";
      when 1848 => r := x"3e8d71543f868db7";
      when 1849 => r := x"3e8d5ec03f8684e1";
      when 1850 => r := x"3e8d4c303f867c0b";
      when 1851 => r := x"3e8d39a33f867337";
      when 1852 => r := x"3e8d271a3f866a64";
      when 1853 => r := x"3e8d14943f866192";
      when 1854 => r := x"3e8d02133f8658c1";
      when 1855 => r := x"3e8cef943f864ff2";
      when 1856 => r := x"3e8cdd1a3f864724";
      when 1857 => r := x"3e8ccaa33f863e56";
      when 1858 => r := x"3e8cb8303f86358a";
      when 1859 => r := x"3e8ca5c03f862cbf";
      when 1860 => r := x"3e8c93543f8623f5";
      when 1861 => r := x"3e8c80ec3f861b2d";
      when 1862 => r := x"3e8c6e873f861265";
      when 1863 => r := x"3e8c5c263f86099f";
      when 1864 => r := x"3e8c49c83f8600da";
      when 1865 => r := x"3e8c376e3f85f816";
      when 1866 => r := x"3e8c25183f85ef53";
      when 1867 => r := x"3e8c12c53f85e691";
      when 1868 => r := x"3e8c00763f85ddd1";
      when 1869 => r := x"3e8bee2a3f85d511";
      when 1870 => r := x"3e8bdbe23f85cc53";
      when 1871 => r := x"3e8bc99e3f85c396";
      when 1872 => r := x"3e8bb75d3f85bada";
      when 1873 => r := x"3e8ba5203f85b21f";
      when 1874 => r := x"3e8b92e63f85a965";
      when 1875 => r := x"3e8b80b03f85a0ac";
      when 1876 => r := x"3e8b6e7d3f8597f5";
      when 1877 => r := x"3e8b5c4e3f858f3f";
      when 1878 => r := x"3e8b4a233f858689";
      when 1879 => r := x"3e8b37fb3f857dd5";
      when 1880 => r := x"3e8b25d73f857522";
      when 1881 => r := x"3e8b13b63f856c71";
      when 1882 => r := x"3e8b01983f8563c0";
      when 1883 => r := x"3e8aef7f3f855b10";
      when 1884 => r := x"3e8add683f855262";
      when 1885 => r := x"3e8acb563f8549b5";
      when 1886 => r := x"3e8ab9473f854109";
      when 1887 => r := x"3e8aa73b3f85385e";
      when 1888 => r := x"3e8a95333f852fb4";
      when 1889 => r := x"3e8a832e3f85270b";
      when 1890 => r := x"3e8a712d3f851e63";
      when 1891 => r := x"3e8a5f303f8515bd";
      when 1892 => r := x"3e8a4d363f850d17";
      when 1893 => r := x"3e8a3b3f3f850473";
      when 1894 => r := x"3e8a294c3f84fbd0";
      when 1895 => r := x"3e8a175d3f84f32e";
      when 1896 => r := x"3e8a05713f84ea8d";
      when 1897 => r := x"3e89f3883f84e1ed";
      when 1898 => r := x"3e89e1a33f84d94f";
      when 1899 => r := x"3e89cfc13f84d0b1";
      when 1900 => r := x"3e89bde33f84c815";
      when 1901 => r := x"3e89ac083f84bf79";
      when 1902 => r := x"3e899a313f84b6df";
      when 1903 => r := x"3e89885e3f84ae46";
      when 1904 => r := x"3e89768d3f84a5ae";
      when 1905 => r := x"3e8964c13f849d17";
      when 1906 => r := x"3e8952f73f849481";
      when 1907 => r := x"3e8941313f848bed";
      when 1908 => r := x"3e892f6f3f848359";
      when 1909 => r := x"3e891db03f847ac7";
      when 1910 => r := x"3e890bf43f847236";
      when 1911 => r := x"3e88fa3c3f8469a5";
      when 1912 => r := x"3e88e8883f846116";
      when 1913 => r := x"3e88d6d63f845888";
      when 1914 => r := x"3e88c5293f844ffb";
      when 1915 => r := x"3e88b37e3f844770";
      when 1916 => r := x"3e88a1d73f843ee5";
      when 1917 => r := x"3e8890343f84365b";
      when 1918 => r := x"3e887e933f842dd3";
      when 1919 => r := x"3e886cf73f84254c";
      when 1920 => r := x"3e885b5d3f841cc5";
      when 1921 => r := x"3e8849c83f841440";
      when 1922 => r := x"3e8838353f840bbc";
      when 1923 => r := x"3e8826a63f840339";
      when 1924 => r := x"3e88151a3f83fab7";
      when 1925 => r := x"3e8803923f83f237";
      when 1926 => r := x"3e87f20d3f83e9b7";
      when 1927 => r := x"3e87e08b3f83e138";
      when 1928 => r := x"3e87cf0d3f83d8bb";
      when 1929 => r := x"3e87bd923f83d03e";
      when 1930 => r := x"3e87ac1b3f83c7c3";
      when 1931 => r := x"3e879aa73f83bf49";
      when 1932 => r := x"3e8789363f83b6d0";
      when 1933 => r := x"3e8777c93f83ae58";
      when 1934 => r := x"3e87665f3f83a5e1";
      when 1935 => r := x"3e8754f83f839d6b";
      when 1936 => r := x"3e8743953f8394f6";
      when 1937 => r := x"3e8732353f838c82";
      when 1938 => r := x"3e8720d93f838410";
      when 1939 => r := x"3e870f803f837b9e";
      when 1940 => r := x"3e86fe2a3f83732e";
      when 1941 => r := x"3e86ecd73f836abf";
      when 1942 => r := x"3e86db883f836250";
      when 1943 => r := x"3e86ca3c3f8359e3";
      when 1944 => r := x"3e86b8f43f835177";
      when 1945 => r := x"3e86a7ae3f83490c";
      when 1946 => r := x"3e86966c3f8340a2";
      when 1947 => r := x"3e86852e3f833839";
      when 1948 => r := x"3e8673f33f832fd1";
      when 1949 => r := x"3e8662bb3f83276b";
      when 1950 => r := x"3e8651863f831f05";
      when 1951 => r := x"3e8640553f8316a1";
      when 1952 => r := x"3e862f273f830e3d";
      when 1953 => r := x"3e861dfc3f8305db";
      when 1954 => r := x"3e860cd43f82fd79";
      when 1955 => r := x"3e85fbb03f82f519";
      when 1956 => r := x"3e85ea8f3f82ecba";
      when 1957 => r := x"3e85d9723f82e45c";
      when 1958 => r := x"3e85c8573f82dbff";
      when 1959 => r := x"3e85b7403f82d3a3";
      when 1960 => r := x"3e85a62d3f82cb48";
      when 1961 => r := x"3e85951c3f82c2ee";
      when 1962 => r := x"3e85840f3f82ba95";
      when 1963 => r := x"3e8573053f82b23d";
      when 1964 => r := x"3e8561fe3f82a9e7";
      when 1965 => r := x"3e8550fb3f82a191";
      when 1966 => r := x"3e853ffb3f82993d";
      when 1967 => r := x"3e852efe3f8290e9";
      when 1968 => r := x"3e851e043f828897";
      when 1969 => r := x"3e850d0e3f828045";
      when 1970 => r := x"3e84fc1a3f8277f5";
      when 1971 => r := x"3e84eb2a3f826fa6";
      when 1972 => r := x"3e84da3e3f826758";
      when 1973 => r := x"3e84c9543f825f0b";
      when 1974 => r := x"3e84b86e3f8256bf";
      when 1975 => r := x"3e84a78b3f824e74";
      when 1976 => r := x"3e8496ab3f82462a";
      when 1977 => r := x"3e8485ce3f823de1";
      when 1978 => r := x"3e8474f53f823599";
      when 1979 => r := x"3e84641f3f822d52";
      when 1980 => r := x"3e84534c3f82250c";
      when 1981 => r := x"3e84427c3f821cc8";
      when 1982 => r := x"3e8431b03f821484";
      when 1983 => r := x"3e8420e63f820c42";
      when 1984 => r := x"3e8410203f820400";
      when 1985 => r := x"3e83ff5d3f81fbbf";
      when 1986 => r := x"3e83ee9d3f81f380";
      when 1987 => r := x"3e83dde13f81eb42";
      when 1988 => r := x"3e83cd273f81e304";
      when 1989 => r := x"3e83bc713f81dac8";
      when 1990 => r := x"3e83abbe3f81d28d";
      when 1991 => r := x"3e839b0e3f81ca53";
      when 1992 => r := x"3e838a613f81c219";
      when 1993 => r := x"3e8379b83f81b9e1";
      when 1994 => r := x"3e8369123f81b1aa";
      when 1995 => r := x"3e83586e3f81a974";
      when 1996 => r := x"3e8347ce3f81a13f";
      when 1997 => r := x"3e8337313f81990b";
      when 1998 => r := x"3e8326983f8190d8";
      when 1999 => r := x"3e8316013f8188a6";
      when 2000 => r := x"3e83056e3f818075";
      when 2001 => r := x"3e82f4dd3f817846";
      when 2002 => r := x"3e82e4503f817017";
      when 2003 => r := x"3e82d3c63f8167e9";
      when 2004 => r := x"3e82c33f3f815fbc";
      when 2005 => r := x"3e82b2bb3f815791";
      when 2006 => r := x"3e82a23b3f814f66";
      when 2007 => r := x"3e8291bd3f81473c";
      when 2008 => r := x"3e8281433f813f14";
      when 2009 => r := x"3e8270cc3f8136ec";
      when 2010 => r := x"3e8260583f812ec6";
      when 2011 => r := x"3e824fe73f8126a0";
      when 2012 => r := x"3e823f793f811e7c";
      when 2013 => r := x"3e822f0e3f811658";
      when 2014 => r := x"3e821ea63f810e36";
      when 2015 => r := x"3e820e413f810614";
      when 2016 => r := x"3e81fde03f80fdf4";
      when 2017 => r := x"3e81ed813f80f5d5";
      when 2018 => r := x"3e81dd263f80edb6";
      when 2019 => r := x"3e81ccce3f80e599";
      when 2020 => r := x"3e81bc793f80dd7d";
      when 2021 => r := x"3e81ac273f80d562";
      when 2022 => r := x"3e819bd83f80cd47";
      when 2023 => r := x"3e818b8c3f80c52e";
      when 2024 => r := x"3e817b433f80bd16";
      when 2025 => r := x"3e816afd3f80b4ff";
      when 2026 => r := x"3e815aba3f80ace8";
      when 2027 => r := x"3e814a7b3f80a4d3";
      when 2028 => r := x"3e813a3e3f809cbf";
      when 2029 => r := x"3e812a053f8094ac";
      when 2030 => r := x"3e8119ce3f808c9a";
      when 2031 => r := x"3e81099b3f808489";
      when 2032 => r := x"3e80f96a3f807c79";
      when 2033 => r := x"3e80e93d3f80746a";
      when 2034 => r := x"3e80d9133f806c5c";
      when 2035 => r := x"3e80c8eb3f80644e";
      when 2036 => r := x"3e80b8c73f805c42";
      when 2037 => r := x"3e80a8a63f805437";
      when 2038 => r := x"3e8098883f804c2d";
      when 2039 => r := x"3e80886d3f804424";
      when 2040 => r := x"3e8078553f803c1c";
      when 2041 => r := x"3e8068403f803415";
      when 2042 => r := x"3e80582e3f802c0f";
      when 2043 => r := x"3e80481f3f80240a";
      when 2044 => r := x"3e8038133f801c06";
      when 2045 => r := x"3e80280a3f801403";
      when 2046 => r := x"3e8018043f800c01";
      when 2047 => r := x"3e8008013f800400";
      when others => r := (others => '0');      -- 0 ~ 2047 まであるのであり得ない。
    end case;
    return r;
  end table;

  component fadd
    port(A : in  std_logic_vector(31 downto 0);
         B : in  std_logic_vector(31 downto 0);
         S : out std_logic_vector(31 downto 0));
  end component;

  component fmul
    port(A : in  std_logic_vector(31 downto 0);
         B : in  std_logic_vector(31 downto 0);
         S : out std_logic_vector(31 downto 0));
  end component; 
  
  constant nan   : std_logic_vector(31 downto 0) := x"7fffffff";
  constant zero  : std_logic_vector(31 downto 0) := x"00000000";
  constant nzero : std_logic_vector(31 downto 0) := x"80000000";
  constant inf   : std_logic_vector(31 downto 0) := x"7f800000";
  constant ninf  : std_logic_vector(31 downto 0) := x"ff800000";

  signal s1,s2,s3,s4,s5 : std_logic_vector(31 downto 0);

begin

  -- Component Instantiation
  fadd_connect : fadd port map(
    A => s3,
    B => s4,
    S => s5);

  fmul_connect : fmul port map(
    A => s1,
    B => s2,
    S => s3);

  do_finv : process(A, s1, s2, s3, s4, s5)
    variable org      : std_logic_vector(31 downto 0);
    variable result   : std_logic_vector(31 downto 0);
    variable fraction : std_logic_vector(31 downto 0);
    variable d        : std_logic_vector(7 downto 0);
    variable index    : std_logic_vector(10 downto 0);
    variable ab_unit  : std_logic_vector(63 downto 0);
    variable ka,kb,temp : std_logic_vector(31 downto 0);   --変更
  begin

    if is_metavalue(A) then
      S <= (others => 'X');
    else
      org := A;

      if (org(30 downto 23) = 255 and org(22 downto 0) /= 0) then
        result := nan;
      elsif org(31) = '0' and org(30 downto 23) = 0 then
        result := inf;
      elsif org(31) = '1' and org(30 downto 23) = 0 then
        result := ninf;
      elsif org = inf then
        result := zero;
      elsif org = ninf then
        result := nzero;
      else
        if org(22 downto 0) = 0 then
          result := org;
          if org(30 downto 23) >= 127 then
            d := org(30 downto 23) - 127;
            result(30 downto 23) := 127 - d;
          else
            d := 127 - org(30 downto 23);
            result(30 downto 23) := 127 + d;
          end if;
        else
          fraction := org;
          fraction(31) := '0';
          fraction(30 downto 23) := "01111111";
          index := fraction(22 downto 12);
          ab_unit := table(index);
          ka := ab_unit(63 downto 32);
          kb := ab_unit(31 downto 0);
          ka(31) := '1';

          s1 <= ka;
          s2 <= fraction;
          s4 <= kb;
          temp := s5;

          result(31) := org(31);
          if org(30 downto 23) >= 127 then
            d := org(30 downto 23) - 127;
            if d < 126 then
              result(30 downto 23) := 126 - d; -- 127 - d - 1
              result(22 downto 0)  := temp(22 downto 0);
            else
              result(30 downto 0) := "000" & x"0000000";
            end if;
          else
            d := 127 - org(30 downto 23);
            result(30 downto 23) := 126 + d; -- 127 + d - 1
            result(22 downto 0)  := temp(22 downto 0);
          end if;
        end if;
      end if;

      S <= result;

    end if;
  end process;
end blackbox;
