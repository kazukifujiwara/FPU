library IEEE;
use IEEE.std_logic_1164.all;

package finv_p is

  component finv is
    port (
      a : in std_logic_vector(31 downto 0);
      s : out std_logic_vector(31 downto 0));
  end component;

end package;


library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_misc.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

library work;
use work.fpu_common_p.all;

entity finv is
  port ( A : in  std_logic_vector(31 downto 0);
         S : out std_logic_vector(31 downto 0));
end entity finv;

architecture blackbox of FINV is

  -- a(32bit) & b(32bit) の計64bitを返す
  function table(index: std_logic_vector(10 downto 0))
    return std_logic_vector
  is
    variable r : std_logic_vector(63 downto 0);
  begin
    case conv_integer(index) is
      when    0 => r := x"3f7fc0103fffe007";
      when    1 => r := x"3f7f40703fffa027";
      when    2 => r := x"3f7ec12f3fff6067";
      when    3 => r := x"3f7e424d3fff20c6";
      when    4 => r := x"3f7dc3ca3ffee146";
      when    5 => r := x"3f7d45a63ffea1e4";
      when    6 => r := x"3f7cc7df3ffe62a3";
      when    7 => r := x"3f7c4a763ffe2380";
      when    8 => r := x"3f7bcd6a3ffde47d";
      when    9 => r := x"3f7b50bb3ffda59a";
      when   10 => r := x"3f7ad4683ffd66d5";
      when   11 => r := x"3f7a58723ffd282f";
      when   12 => r := x"3f79dcd83ffce9a9";
      when   13 => r := x"3f7961993ffcab41";
      when   14 => r := x"3f78e6b53ffc6cf8";
      when   15 => r := x"3f786c2b3ffc2ece";
      when   16 => r := x"3f77f1fd3ffbf0c2";
      when   17 => r := x"3f7778283ffbb2d5";
      when   18 => r := x"3f76fead3ffb7506";
      when   19 => r := x"3f76858b3ffb3755";
      when   20 => r := x"3f760cc23ffaf9c3";
      when   21 => r := x"3f7594523ffabc4f";
      when   22 => r := x"3f751c3b3ffa7ef9";
      when   23 => r := x"3f74a47b3ffa41c1";
      when   24 => r := x"3f742d133ffa04a6";
      when   25 => r := x"3f73b6033ff9c7aa";
      when   26 => r := x"3f733f493ff98acb";
      when   27 => r := x"3f72c8e63ff94e0a";
      when   28 => r := x"3f7252d93ff91167";
      when   29 => r := x"3f71dd233ff8d4e1";
      when   30 => r := x"3f7167c23ff89878";
      when   31 => r := x"3f70f2b63ff85c2d";
      when   32 => r := x"3f707e003ff81fff";
      when   33 => r := x"3f70099e3ff7e3ee";
      when   34 => r := x"3f6f95913ff7a7fa";
      when   35 => r := x"3f6f21d83ff76c23";
      when   36 => r := x"3f6eae723ff73069";
      when   37 => r := x"3f6e3b603ff6f4cc";
      when   38 => r := x"3f6dc8a13ff6b94b";
      when   39 => r := x"3f6d56353ff67de7";
      when   40 => r := x"3f6ce41b3ff642a0";
      when   41 => r := x"3f6c72543ff60775";
      when   42 => r := x"3f6c00df3ff5cc67";
      when   43 => r := x"3f6b8fbb3ff59175";
      when   44 => r := x"3f6b1ee83ff5569f";
      when   45 => r := x"3f6aae673ff51be5";
      when   46 => r := x"3f6a3e363ff4e148";
      when   47 => r := x"3f69ce553ff4a6c6";
      when   48 => r := x"3f695ec43ff46c61";
      when   49 => r := x"3f68ef843ff43217";
      when   50 => r := x"3f6880933ff3f7e9";
      when   51 => r := x"3f6811f03ff3bdd7";
      when   52 => r := x"3f67a39d3ff383e0";
      when   53 => r := x"3f6735993ff34a05";
      when   54 => r := x"3f66c7e23ff31045";
      when   55 => r := x"3f665a7a3ff2d6a1";
      when   56 => r := x"3f65ed603ff29d18";
      when   57 => r := x"3f6580933ff263aa";
      when   58 => r := x"3f6514133ff22a57";
      when   59 => r := x"3f64a7e03ff1f120";
      when   60 => r := x"3f643bf93ff1b803";
      when   61 => r := x"3f63d05f3ff17f02";
      when   62 => r := x"3f6365113ff1461b";
      when   63 => r := x"3f62fa0f3ff10d4f";
      when   64 => r := x"3f628f583ff0d49e";
      when   65 => r := x"3f6224ec3ff09c08";
      when   66 => r := x"3f61bacb3ff0638c";
      when   67 => r := x"3f6150f53ff02b2a";
      when   68 => r := x"3f60e7693feff2e3";
      when   69 => r := x"3f607e273fefbab6";
      when   70 => r := x"3f6015303fef82a4";
      when   71 => r := x"3f5fac813fef4aac";
      when   72 => r := x"3f5f441c3fef12ce";
      when   73 => r := x"3f5edc003feedb0a";
      when   74 => r := x"3f5e742d3feea360";
      when   75 => r := x"3f5e0ca23fee6bd0";
      when   76 => r := x"3f5da55f3fee3459";
      when   77 => r := x"3f5d3e653fedfcfd";
      when   78 => r := x"3f5cd7b23fedc5ba";
      when   79 => r := x"3f5c71473fed8e91";
      when   80 => r := x"3f5c0b223fed5782";
      when   81 => r := x"3f5ba5453fed208b";
      when   82 => r := x"3f5b3fae3fece9af";
      when   83 => r := x"3f5ada5e3fecb2ec";
      when   84 => r := x"3f5a75543fec7c42";
      when   85 => r := x"3f5a10903fec45b1";
      when   86 => r := x"3f59ac113fec0f39";
      when   87 => r := x"3f5947d83febd8db";
      when   88 => r := x"3f58e3e43feba295";
      when   89 => r := x"3f5880353feb6c69";
      when   90 => r := x"3f581ccb3feb3655";
      when   91 => r := x"3f57b9a53feb005a";
      when   92 => r := x"3f5756c33feaca78";
      when   93 => r := x"3f56f4253fea94af";
      when   94 => r := x"3f5691cb3fea5efe";
      when   95 => r := x"3f562fb43fea2966";
      when   96 => r := x"3f55cde03fe9f3e6";
      when   97 => r := x"3f556c503fe9be7f";
      when   98 => r := x"3f550b023fe98930";
      when   99 => r := x"3f54a9f73fe953fa";
      when  100 => r := x"3f54492d3fe91edb";
      when  101 => r := x"3f53e8a63fe8e9d5";
      when  102 => r := x"3f5388613fe8b4e7";
      when  103 => r := x"3f53285d3fe88011";
      when  104 => r := x"3f52c89b3fe84b53";
      when  105 => r := x"3f5269193fe816ac";
      when  106 => r := x"3f5209d93fe7e21e";
      when  107 => r := x"3f51aad93fe7ada7";
      when  108 => r := x"3f514c193fe77949";
      when  109 => r := x"3f50ed9a3fe74501";
      when  110 => r := x"3f508f5a3fe710d2";
      when  111 => r := x"3f50315b3fe6dcba";
      when  112 => r := x"3f4fd39a3fe6a8b9";
      when  113 => r := x"3f4f761a3fe674d0";
      when  114 => r := x"3f4f18d83fe640fe";
      when  115 => r := x"3f4ebbd53fe60d43";
      when  116 => r := x"3f4e5f103fe5d9a0";
      when  117 => r := x"3f4e028a3fe5a614";
      when  118 => r := x"3f4da6423fe5729f";
      when  119 => r := x"3f4d4a383fe53f41";
      when  120 => r := x"3f4cee6c3fe50bfa";
      when  121 => r := x"3f4c92dd3fe4d8c9";
      when  122 => r := x"3f4c378c3fe4a5b0";
      when  123 => r := x"3f4bdc773fe472ae";
      when  124 => r := x"3f4b81a03fe43fc2";
      when  125 => r := x"3f4b27053fe40ced";
      when  126 => r := x"3f4acca73fe3da2e";
      when  127 => r := x"3f4a72853fe3a787";
      when  128 => r := x"3f4a189f3fe374f5";
      when  129 => r := x"3f49bef53fe3427a";
      when  130 => r := x"3f4965863fe31016";
      when  131 => r := x"3f490c533fe2ddc7";
      when  132 => r := x"3f48b35b3fe2ab8f";
      when  133 => r := x"3f485a9e3fe2796e";
      when  134 => r := x"3f48021c3fe24762";
      when  135 => r := x"3f47a9d43fe2156d";
      when  136 => r := x"3f4751c73fe1e38d";
      when  137 => r := x"3f46f9f43fe1b1c4";
      when  138 => r := x"3f46a25b3fe18010";
      when  139 => r := x"3f464afc3fe14e72";
      when  140 => r := x"3f45f3d73fe11ceb";
      when  141 => r := x"3f459cea3fe0eb79";
      when  142 => r := x"3f4546373fe0ba1c";
      when  143 => r := x"3f44efbd3fe088d5";
      when  144 => r := x"3f44997c3fe057a4";
      when  145 => r := x"3f4443743fe02689";
      when  146 => r := x"3f43eda43fdff583";
      when  147 => r := x"3f43980c3fdfc492";
      when  148 => r := x"3f4342ac3fdf93b6";
      when  149 => r := x"3f42ed843fdf62f0";
      when  150 => r := x"3f4298943fdf3240";
      when  151 => r := x"3f4243db3fdf01a4";
      when  152 => r := x"3f41ef593fded11e";
      when  153 => r := x"3f419b0f3fdea0ac";
      when  154 => r := x"3f4146fb3fde7050";
      when  155 => r := x"3f40f31e3fde4009";
      when  156 => r := x"3f409f783fde0fd7";
      when  157 => r := x"3f404c083fdddfb9";
      when  158 => r := x"3f3ff8ce3fddafb1";
      when  159 => r := x"3f3fa5ca3fdd7fbd";
      when  160 => r := x"3f3f52fc3fdd4fde";
      when  161 => r := x"3f3f00643fdd2013";
      when  162 => r := x"3f3eae013fdcf05d";
      when  163 => r := x"3f3e5bd33fdcc0bc";
      when  164 => r := x"3f3e09db3fdc912f";
      when  165 => r := x"3f3db8173fdc61b7";
      when  166 => r := x"3f3d66883fdc3253";
      when  167 => r := x"3f3d152e3fdc0304";
      when  168 => r := x"3f3cc4083fdbd3c9";
      when  169 => r := x"3f3c73163fdba4a2";
      when  170 => r := x"3f3c22583fdb758f";
      when  171 => r := x"3f3bd1ce3fdb4691";
      when  172 => r := x"3f3b81783fdb17a6";
      when  173 => r := x"3f3b31553fdae8d0";
      when  174 => r := x"3f3ae1653fdaba0e";
      when  175 => r := x"3f3a91a93fda8b5f";
      when  176 => r := x"3f3a42203fda5cc5";
      when  177 => r := x"3f39f2c93fda2e3e";
      when  178 => r := x"3f39a3a53fd9ffcb";
      when  179 => r := x"3f3954b43fd9d16c";
      when  180 => r := x"3f3905f53fd9a321";
      when  181 => r := x"3f38b7683fd974e9";
      when  182 => r := x"3f38690d3fd946c5";
      when  183 => r := x"3f381ae43fd918b5";
      when  184 => r := x"3f37ccec3fd8eab8";
      when  185 => r := x"3f377f263fd8bcce";
      when  186 => r := x"3f3731923fd88ef8";
      when  187 => r := x"3f36e42e3fd86135";
      when  188 => r := x"3f3696fc3fd83386";
      when  189 => r := x"3f3649fa3fd805ea";
      when  190 => r := x"3f35fd293fd7d861";
      when  191 => r := x"3f35b0883fd7aaeb";
      when  192 => r := x"3f3564183fd77d89";
      when  193 => r := x"3f3517d83fd75039";
      when  194 => r := x"3f34cbc83fd722fd";
      when  195 => r := x"3f347fe83fd6f5d3";
      when  196 => r := x"3f3434383fd6c8bd";
      when  197 => r := x"3f33e8b73fd69bb9";
      when  198 => r := x"3f339d663fd66ec8";
      when  199 => r := x"3f3352443fd641eb";
      when  200 => r := x"3f3307513fd6151f";
      when  201 => r := x"3f32bc8d3fd5e867";
      when  202 => r := x"3f3271f83fd5bbc1";
      when  203 => r := x"3f3227913fd58f2e";
      when  204 => r := x"3f31dd593fd562ad";
      when  205 => r := x"3f3193503fd5363f";
      when  206 => r := x"3f3149743fd509e4";
      when  207 => r := x"3f30ffc73fd4dd9a";
      when  208 => r := x"3f30b6473fd4b164";
      when  209 => r := x"3f306cf53fd4853f";
      when  210 => r := x"3f3023d13fd4592d";
      when  211 => r := x"3f2fdada3fd42d2d";
      when  212 => r := x"3f2f92113fd40140";
      when  213 => r := x"3f2f49743fd3d564";
      when  214 => r := x"3f2f01053fd3a99b";
      when  215 => r := x"3f2eb8c23fd37de4";
      when  216 => r := x"3f2e70ad3fd3523f";
      when  217 => r := x"3f2e28c33fd326ab";
      when  218 => r := x"3f2de1073fd2fb2a";
      when  219 => r := x"3f2d99763fd2cfbb";
      when  220 => r := x"3f2d52123fd2a45d";
      when  221 => r := x"3f2d0ada3fd27912";
      when  222 => r := x"3f2cc3cd3fd24dd8";
      when  223 => r := x"3f2c7cec3fd222b0";
      when  224 => r := x"3f2c36373fd1f799";
      when  225 => r := x"3f2befad3fd1cc95";
      when  226 => r := x"3f2ba94f3fd1a1a2";
      when  227 => r := x"3f2b631c3fd176c0";
      when  228 => r := x"3f2b1d143fd14bf0";
      when  229 => r := x"3f2ad7363fd12132";
      when  230 => r := x"3f2a91843fd0f684";
      when  231 => r := x"3f2a4bfc3fd0cbe9";
      when  232 => r := x"3f2a069e3fd0a15e";
      when  233 => r := x"3f29c16b3fd076e5";
      when  234 => r := x"3f297c623fd04c7e";
      when  235 => r := x"3f2937833fd02227";
      when  236 => r := x"3f28f2cf3fcff7e2";
      when  237 => r := x"3f28ae433fcfcdae";
      when  238 => r := x"3f2869e23fcfa38b";
      when  239 => r := x"3f2825aa3fcf7979";
      when  240 => r := x"3f27e19c3fcf4f78";
      when  241 => r := x"3f279db73fcf2588";
      when  242 => r := x"3f2759fb3fcefba9";
      when  243 => r := x"3f2716683fced1db";
      when  244 => r := x"3f26d2fe3fcea81e";
      when  245 => r := x"3f268fbc3fce7e71";
      when  246 => r := x"3f264ca43fce54d6";
      when  247 => r := x"3f2609b33fce2b4b";
      when  248 => r := x"3f25c6ec3fce01d1";
      when  249 => r := x"3f25844c3fcdd868";
      when  250 => r := x"3f2541d53fcdaf0f";
      when  251 => r := x"3f24ff853fcd85c7";
      when  252 => r := x"3f24bd5e3fcd5c8f";
      when  253 => r := x"3f247b5e3fcd3368";
      when  254 => r := x"3f2439863fcd0a51";
      when  255 => r := x"3f23f7d53fcce14b";
      when  256 => r := x"3f23b64c3fccb856";
      when  257 => r := x"3f2374ea3fcc8f70";
      when  258 => r := x"3f2333af3fcc669b";
      when  259 => r := x"3f22f29c3fcc3dd6";
      when  260 => r := x"3f22b1af3fcc1522";
      when  261 => r := x"3f2270e93fcbec7d";
      when  262 => r := x"3f2230493fcbc3e9";
      when  263 => r := x"3f21efd03fcb9b65";
      when  264 => r := x"3f21af7e3fcb72f1";
      when  265 => r := x"3f216f513fcb4a8d";
      when  266 => r := x"3f212f4b3fcb223a";
      when  267 => r := x"3f20ef6b3fcaf9f6";
      when  268 => r := x"3f20afb13fcad1c2";
      when  269 => r := x"3f20701d3fcaa99e";
      when  270 => r := x"3f2030ae3fca818a";
      when  271 => r := x"3f1ff1653fca5986";
      when  272 => r := x"3f1fb2423fca3191";
      when  273 => r := x"3f1f73443fca09ac";
      when  274 => r := x"3f1f346b3fc9e1d7";
      when  275 => r := x"3f1ef5b73fc9ba12";
      when  276 => r := x"3f1eb7283fc9925d";
      when  277 => r := x"3f1e78be3fc96ab7";
      when  278 => r := x"3f1e3a793fc94320";
      when  279 => r := x"3f1dfc593fc91b99";
      when  280 => r := x"3f1dbe5d3fc8f422";
      when  281 => r := x"3f1d80863fc8ccba";
      when  282 => r := x"3f1d42d33fc8a562";
      when  283 => r := x"3f1d05443fc87e19";
      when  284 => r := x"3f1cc7d93fc856df";
      when  285 => r := x"3f1c8a933fc82fb5";
      when  286 => r := x"3f1c4d703fc8089a";
      when  287 => r := x"3f1c10713fc7e18e";
      when  288 => r := x"3f1bd3963fc7ba92";
      when  289 => r := x"3f1b96de3fc793a4";
      when  290 => r := x"3f1b5a493fc76cc6";
      when  291 => r := x"3f1b1dd93fc745f7";
      when  292 => r := x"3f1ae18b3fc71f37";
      when  293 => r := x"3f1aa5603fc6f886";
      when  294 => r := x"3f1a69593fc6d1e4";
      when  295 => r := x"3f1a2d743fc6ab52";
      when  296 => r := x"3f19f1b23fc684ce";
      when  297 => r := x"3f19b6133fc65e59";
      when  298 => r := x"3f197a973fc637f3";
      when  299 => r := x"3f193f3d3fc6119b";
      when  300 => r := x"3f1904053fc5eb53";
      when  301 => r := x"3f18c8f03fc5c519";
      when  302 => r := x"3f188dfd3fc59eef";
      when  303 => r := x"3f18532c3fc578d2";
      when  304 => r := x"3f18187d3fc552c5";
      when  305 => r := x"3f17ddf03fc52cc6";
      when  306 => r := x"3f17a3853fc506d6";
      when  307 => r := x"3f17693b3fc4e0f4";
      when  308 => r := x"3f172f133fc4bb21";
      when  309 => r := x"3f16f50d3fc4955d";
      when  310 => r := x"3f16bb273fc46fa7";
      when  311 => r := x"3f1681643fc449ff";
      when  312 => r := x"3f1647c13fc42466";
      when  313 => r := x"3f160e3f3fc3fedb";
      when  314 => r := x"3f15d4df3fc3d95f";
      when  315 => r := x"3f159b9f3fc3b3f1";
      when  316 => r := x"3f1562803fc38e91";
      when  317 => r := x"3f1529823fc36940";
      when  318 => r := x"3f14f0a43fc343fc";
      when  319 => r := x"3f14b7e73fc31ec7";
      when  320 => r := x"3f147f4a3fc2f9a0";
      when  321 => r := x"3f1446cd3fc2d488";
      when  322 => r := x"3f140e713fc2af7d";
      when  323 => r := x"3f13d6353fc28a80";
      when  324 => r := x"3f139e193fc26592";
      when  325 => r := x"3f13661c3fc240b1";
      when  326 => r := x"3f132e403fc21bdf";
      when  327 => r := x"3f12f6833fc1f71a";
      when  328 => r := x"3f12bee63fc1d264";
      when  329 => r := x"3f1287693fc1adbb";
      when  330 => r := x"3f12500b3fc18920";
      when  331 => r := x"3f1218cc3fc16493";
      when  332 => r := x"3f11e1ad3fc14013";
      when  333 => r := x"3f11aaac3fc11ba2";
      when  334 => r := x"3f1173cb3fc0f73e";
      when  335 => r := x"3f113d093fc0d2e8";
      when  336 => r := x"3f1106663fc0aea0";
      when  337 => r := x"3f10cfe13fc08a65";
      when  338 => r := x"3f10997c3fc06638";
      when  339 => r := x"3f1063343fc04218";
      when  340 => r := x"3f102d0c3fc01e06";
      when  341 => r := x"3f0ff7023fbffa01";
      when  342 => r := x"3f0fc1163fbfd60a";
      when  343 => r := x"3f0f8b483fbfb221";
      when  344 => r := x"3f0f55993fbf8e45";
      when  345 => r := x"3f0f20083fbf6a76";
      when  346 => r := x"3f0eea953fbf46b5";
      when  347 => r := x"3f0eb53f3fbf2301";
      when  348 => r := x"3f0e80083fbeff5a";
      when  349 => r := x"3f0e4aee3fbedbc1";
      when  350 => r := x"3f0e15f23fbeb835";
      when  351 => r := x"3f0de1143fbe94b6";
      when  352 => r := x"3f0dac533fbe7144";
      when  353 => r := x"3f0d77af3fbe4de0";
      when  354 => r := x"3f0d43293fbe2a88";
      when  355 => r := x"3f0d0ec03fbe073e";
      when  356 => r := x"3f0cda743fbde401";
      when  357 => r := x"3f0ca6453fbdc0d1";
      when  358 => r := x"3f0c72333fbd9dae";
      when  359 => r := x"3f0c3e3e3fbd7a98";
      when  360 => r := x"3f0c0a663fbd578f";
      when  361 => r := x"3f0bd6aa3fbd3492";
      when  362 => r := x"3f0ba30c3fbd11a3";
      when  363 => r := x"3f0b6f893fbceec1";
      when  364 => r := x"3f0b3c243fbccbeb";
      when  365 => r := x"3f0b08da3fbca923";
      when  366 => r := x"3f0ad5ad3fbc8667";
      when  367 => r := x"3f0aa29c3fbc63b8";
      when  368 => r := x"3f0a6fa83fbc4116";
      when  369 => r := x"3f0a3ccf3fbc1e80";
      when  370 => r := x"3f0a0a133fbbfbf7";
      when  371 => r := x"3f09d7723fbbd97b";
      when  372 => r := x"3f09a4ed3fbbb70c";
      when  373 => r := x"3f0972843fbb94a9";
      when  374 => r := x"3f0940373fbb7252";
      when  375 => r := x"3f090e053fbb5008";
      when  376 => r := x"3f08dbef3fbb2dcb";
      when  377 => r := x"3f08a9f43fbb0b9b";
      when  378 => r := x"3f0878143fbae976";
      when  379 => r := x"3f0846503fbac75e";
      when  380 => r := x"3f0814a73fbaa553";
      when  381 => r := x"3f07e3193fba8354";
      when  382 => r := x"3f07b1a63fba6162";
      when  383 => r := x"3f07804e3fba3f7b";
      when  384 => r := x"3f074f113fba1da1";
      when  385 => r := x"3f071def3fb9fbd4";
      when  386 => r := x"3f06ece83fb9da12";
      when  387 => r := x"3f06bbfb3fb9b85d";
      when  388 => r := x"3f068b293fb996b4";
      when  389 => r := x"3f065a713fb97518";
      when  390 => r := x"3f0629d43fb95387";
      when  391 => r := x"3f05f9513fb93203";
      when  392 => r := x"3f05c8e93fb9108a";
      when  393 => r := x"3f05989a3fb8ef1e";
      when  394 => r := x"3f0568663fb8cdbe";
      when  395 => r := x"3f05384c3fb8ac6a";
      when  396 => r := x"3f05084c3fb88b22";
      when  397 => r := x"3f04d8663fb869e6";
      when  398 => r := x"3f04a8993fb848b6";
      when  399 => r := x"3f0478e73fb82792";
      when  400 => r := x"3f04494e3fb80679";
      when  401 => r := x"3f0419cf3fb7e56d";
      when  402 => r := x"3f03ea693fb7c46c";
      when  403 => r := x"3f03bb1d3fb7a378";
      when  404 => r := x"3f038bea3fb7828f";
      when  405 => r := x"3f035cd13fb761b2";
      when  406 => r := x"3f032dd13fb740e0";
      when  407 => r := x"3f02feea3fb7201b";
      when  408 => r := x"3f02d01c3fb6ff61";
      when  409 => r := x"3f02a1673fb6deb3";
      when  410 => r := x"3f0272cc3fb6be10";
      when  411 => r := x"3f0244493fb69d79";
      when  412 => r := x"3f0215df3fb67cee";
      when  413 => r := x"3f01e78e3fb65c6e";
      when  414 => r := x"3f01b9553fb63bfa";
      when  415 => r := x"3f018b363fb61b92";
      when  416 => r := x"3f015d2f3fb5fb35";
      when  417 => r := x"3f012f403fb5dae3";
      when  418 => r := x"3f01016a3fb5ba9d";
      when  419 => r := x"3f00d3ac3fb59a62";
      when  420 => r := x"3f00a6063fb57a33";
      when  421 => r := x"3f0078793fb55a0f";
      when  422 => r := x"3f004b043fb539f7";
      when  423 => r := x"3f001da73fb519ea";
      when  424 => r := x"3effe0c43fb4f9e8";
      when  425 => r := x"3eff866a3fb4d9f2";
      when  426 => r := x"3eff2c403fb4ba07";
      when  427 => r := x"3efed2453fb49a27";
      when  428 => r := x"3efe787a3fb47a52";
      when  429 => r := x"3efe1edf3fb45a88";
      when  430 => r := x"3efdc5733fb43aca";
      when  431 => r := x"3efd6c363fb41b17";
      when  432 => r := x"3efd13283fb3fb6f";
      when  433 => r := x"3efcba493fb3dbd2";
      when  434 => r := x"3efc61993fb3bc41";
      when  435 => r := x"3efc09173fb39cba";
      when  436 => r := x"3efbb0c43fb37d3e";
      when  437 => r := x"3efb589f3fb35dce";
      when  438 => r := x"3efb00a93fb33e68";
      when  439 => r := x"3efaa8e03fb31f0e";
      when  440 => r := x"3efa51463fb2ffbe";
      when  441 => r := x"3ef9f9da3fb2e079";
      when  442 => r := x"3ef9a29b3fb2c13f";
      when  443 => r := x"3ef94b8a3fb2a211";
      when  444 => r := x"3ef8f4a73fb282ed";
      when  445 => r := x"3ef89df13fb263d3";
      when  446 => r := x"3ef847683fb244c5";
      when  447 => r := x"3ef7f10c3fb225c2";
      when  448 => r := x"3ef79ade3fb206c9";
      when  449 => r := x"3ef744dc3fb1e7db";
      when  450 => r := x"3ef6ef073fb1c8f8";
      when  451 => r := x"3ef6995f3fb1aa1f";
      when  452 => r := x"3ef643e33fb18b51";
      when  453 => r := x"3ef5ee943fb16c8e";
      when  454 => r := x"3ef599713fb14dd6";
      when  455 => r := x"3ef5447a3fb12f28";
      when  456 => r := x"3ef4efaf3fb11084";
      when  457 => r := x"3ef49b113fb0f1ec";
      when  458 => r := x"3ef4469e3fb0d35e";
      when  459 => r := x"3ef3f2563fb0b4da";
      when  460 => r := x"3ef39e3b3fb09661";
      when  461 => r := x"3ef34a4a3fb077f3";
      when  462 => r := x"3ef2f6863fb0598e";
      when  463 => r := x"3ef2a2ec3fb03b35";
      when  464 => r := x"3ef24f7d3fb01ce6";
      when  465 => r := x"3ef1fc3a3faffea1";
      when  466 => r := x"3ef1a9213fafe067";
      when  467 => r := x"3ef156333fafc237";
      when  468 => r := x"3ef103703fafa411";
      when  469 => r := x"3ef0b0d73faf85f6";
      when  470 => r := x"3ef05e693faf67e5";
      when  471 => r := x"3ef00c253faf49de";
      when  472 => r := x"3eefba0c3faf2be2";
      when  473 => r := x"3eef681c3faf0df0";
      when  474 => r := x"3eef16563faef008";
      when  475 => r := x"3eeec4bb3faed22a";
      when  476 => r := x"3eee73493faeb457";
      when  477 => r := x"3eee22003fae968d";
      when  478 => r := x"3eedd0e13fae78ce";
      when  479 => r := x"3eed7fec3fae5b19";
      when  480 => r := x"3eed2f203fae3d6e";
      when  481 => r := x"3eecde7d3fae1fcd";
      when  482 => r := x"3eec8e033fae0236";
      when  483 => r := x"3eec3db23fade4aa";
      when  484 => r := x"3eebed8b3fadc727";
      when  485 => r := x"3eeb9d8b3fada9ae";
      when  486 => r := x"3eeb4db53fad8c40";
      when  487 => r := x"3eeafe073fad6edb";
      when  488 => r := x"3eeaae813fad5180";
      when  489 => r := x"3eea5f243fad342f";
      when  490 => r := x"3eea0fef3fad16e8";
      when  491 => r := x"3ee9c0e23facf9ab";
      when  492 => r := x"3ee971fe3facdc78";
      when  493 => r := x"3ee923413facbf4f";
      when  494 => r := x"3ee8d4ac3faca22f";
      when  495 => r := x"3ee8863e3fac851a";
      when  496 => r := x"3ee837f93fac680e";
      when  497 => r := x"3ee7e9da3fac4b0c";
      when  498 => r := x"3ee79be33fac2e13";
      when  499 => r := x"3ee74e143fac1125";
      when  500 => r := x"3ee7006b3fabf440";
      when  501 => r := x"3ee6b2ea3fabd765";
      when  502 => r := x"3ee665903fabba93";
      when  503 => r := x"3ee6185c3fab9dcb";
      when  504 => r := x"3ee5cb503fab810d";
      when  505 => r := x"3ee57e6a3fab6458";
      when  506 => r := x"3ee531aa3fab47ad";
      when  507 => r := x"3ee4e5113fab2b0c";
      when  508 => r := x"3ee4989f3fab0e74";
      when  509 => r := x"3ee44c523faaf1e6";
      when  510 => r := x"3ee4002c3faad561";
      when  511 => r := x"3ee3b42c3faab8e6";
      when  512 => r := x"3ee368523faa9c74";
      when  513 => r := x"3ee31c9e3faa800c";
      when  514 => r := x"3ee2d1103faa63ad";
      when  515 => r := x"3ee285a73faa4757";
      when  516 => r := x"3ee23a643faa2b0b";
      when  517 => r := x"3ee1ef463faa0ec9";
      when  518 => r := x"3ee1a44e3fa9f28f";
      when  519 => r := x"3ee1597b3fa9d660";
      when  520 => r := x"3ee10ecd3fa9ba39";
      when  521 => r := x"3ee0c4443fa99e1c";
      when  522 => r := x"3ee079e03fa98208";
      when  523 => r := x"3ee02fa23fa965fd";
      when  524 => r := x"3edfe5883fa949fc";
      when  525 => r := x"3edf9b923fa92e04";
      when  526 => r := x"3edf51c23fa91215";
      when  527 => r := x"3edf08163fa8f630";
      when  528 => r := x"3edebe8e3fa8da53";
      when  529 => r := x"3ede752b3fa8be80";
      when  530 => r := x"3ede2beb3fa8a2b6";
      when  531 => r := x"3edde2d03fa886f5";
      when  532 => r := x"3edd99da3fa86b3d";
      when  533 => r := x"3edd51073fa84f8e";
      when  534 => r := x"3edd08583fa833e9";
      when  535 => r := x"3edcbfcc3fa8184c";
      when  536 => r := x"3edc77653fa7fcb9";
      when  537 => r := x"3edc2f213fa7e12f";
      when  538 => r := x"3edbe7003fa7c5ad";
      when  539 => r := x"3edb9f033fa7aa35";
      when  540 => r := x"3edb572a3fa78ec5";
      when  541 => r := x"3edb0f733fa7735f";
      when  542 => r := x"3edac7e03fa75801";
      when  543 => r := x"3eda806f3fa73cad";
      when  544 => r := x"3eda39223fa72161";
      when  545 => r := x"3ed9f1f83fa7061f";
      when  546 => r := x"3ed9aaf03fa6eae5";
      when  547 => r := x"3ed9640b3fa6cfb4";
      when  548 => r := x"3ed91d493fa6b48c";
      when  549 => r := x"3ed8d6a93fa6996d";
      when  550 => r := x"3ed8902c3fa67e56";
      when  551 => r := x"3ed849d13fa66349";
      when  552 => r := x"3ed803983fa64844";
      when  553 => r := x"3ed7bd813fa62d48";
      when  554 => r := x"3ed7778d3fa61254";
      when  555 => r := x"3ed731ba3fa5f76a";
      when  556 => r := x"3ed6ec0a3fa5dc88";
      when  557 => r := x"3ed6a67b3fa5c1af";
      when  558 => r := x"3ed6610e3fa5a6de";
      when  559 => r := x"3ed61bc33fa58c16";
      when  560 => r := x"3ed5d6993fa57157";
      when  561 => r := x"3ed591913fa556a1";
      when  562 => r := x"3ed54caa3fa53bf3";
      when  563 => r := x"3ed507e43fa5214e";
      when  564 => r := x"3ed4c3403fa506b1";
      when  565 => r := x"3ed47ebd3fa4ec1d";
      when  566 => r := x"3ed43a5b3fa4d191";
      when  567 => r := x"3ed3f61a3fa4b70e";
      when  568 => r := x"3ed3b1f93fa49c94";
      when  569 => r := x"3ed36dfa3fa48222";
      when  570 => r := x"3ed32a1b3fa467b8";
      when  571 => r := x"3ed2e65d3fa44d57";
      when  572 => r := x"3ed2a2c03fa432ff";
      when  573 => r := x"3ed25f433fa418af";
      when  574 => r := x"3ed21be73fa3fe67";
      when  575 => r := x"3ed1d8ab3fa3e428";
      when  576 => r := x"3ed1958f3fa3c9f1";
      when  577 => r := x"3ed152933fa3afc2";
      when  578 => r := x"3ed10fb73fa3959c";
      when  579 => r := x"3ed0ccfc3fa37b7e";
      when  580 => r := x"3ed08a603fa36169";
      when  581 => r := x"3ed047e43fa3475c";
      when  582 => r := x"3ed005883fa32d57";
      when  583 => r := x"3ecfc34c3fa3135a";
      when  584 => r := x"3ecf812f3fa2f966";
      when  585 => r := x"3ecf3f323fa2df7a";
      when  586 => r := x"3ecefd543fa2c596";
      when  587 => r := x"3ecebb963fa2abbb";
      when  588 => r := x"3ece79f73fa291e7";
      when  589 => r := x"3ece38773fa2781c";
      when  590 => r := x"3ecdf7163fa25e59";
      when  591 => r := x"3ecdb5d53fa2449e";
      when  592 => r := x"3ecd74b23fa22aec";
      when  593 => r := x"3ecd33ae3fa21141";
      when  594 => r := x"3eccf2ca3fa1f79f";
      when  595 => r := x"3eccb2043fa1de04";
      when  596 => r := x"3ecc715c3fa1c472";
      when  597 => r := x"3ecc30d33fa1aae8";
      when  598 => r := x"3ecbf0693fa19166";
      when  599 => r := x"3ecbb01d3fa177ec";
      when  600 => r := x"3ecb6ff03fa15e7a";
      when  601 => r := x"3ecb2fe13fa14510";
      when  602 => r := x"3ecaeff03fa12bae";
      when  603 => r := x"3ecab01d3fa11254";
      when  604 => r := x"3eca70693fa0f902";
      when  605 => r := x"3eca30d23fa0dfb8";
      when  606 => r := x"3ec9f1593fa0c676";
      when  607 => r := x"3ec9b1ff3fa0ad3c";
      when  608 => r := x"3ec972c23fa09409";
      when  609 => r := x"3ec933a23fa07adf";
      when  610 => r := x"3ec8f4a13fa061bc";
      when  611 => r := x"3ec8b5bd3fa048a2";
      when  612 => r := x"3ec876f63fa02f8f";
      when  613 => r := x"3ec8384d3fa01684";
      when  614 => r := x"3ec7f9c13f9ffd81";
      when  615 => r := x"3ec7bb533f9fe485";
      when  616 => r := x"3ec77d023f9fcb92";
      when  617 => r := x"3ec73ece3f9fb2a6";
      when  618 => r := x"3ec700b73f9f99c2";
      when  619 => r := x"3ec6c2bd3f9f80e6";
      when  620 => r := x"3ec684e03f9f6812";
      when  621 => r := x"3ec6471f3f9f4f45";
      when  622 => r := x"3ec6097c3f9f3680";
      when  623 => r := x"3ec5cbf53f9f1dc2";
      when  624 => r := x"3ec58e8b3f9f050d";
      when  625 => r := x"3ec5513e3f9eec5f";
      when  626 => r := x"3ec5140d3f9ed3b8";
      when  627 => r := x"3ec4d6f83f9ebb1a";
      when  628 => r := x"3ec49a003f9ea283";
      when  629 => r := x"3ec45d253f9e89f3";
      when  630 => r := x"3ec420653f9e716b";
      when  631 => r := x"3ec3e3c23f9e58eb";
      when  632 => r := x"3ec3a73a3f9e4072";
      when  633 => r := x"3ec36acf3f9e2801";
      when  634 => r := x"3ec32e803f9e0f98";
      when  635 => r := x"3ec2f24d3f9df736";
      when  636 => r := x"3ec2b6353f9ddedb";
      when  637 => r := x"3ec27a393f9dc688";
      when  638 => r := x"3ec23e593f9dae3d";
      when  639 => r := x"3ec202953f9d95f9";
      when  640 => r := x"3ec1c6ec3f9d7dbc";
      when  641 => r := x"3ec18b5f3f9d6587";
      when  642 => r := x"3ec14fed3f9d4d59";
      when  643 => r := x"3ec114963f9d3533";
      when  644 => r := x"3ec0d95b3f9d1d14";
      when  645 => r := x"3ec09e3b3f9d04fc";
      when  646 => r := x"3ec063363f9cecec";
      when  647 => r := x"3ec0284c3f9cd4e4";
      when  648 => r := x"3ebfed7e3f9cbce2";
      when  649 => r := x"3ebfb2ca3f9ca4e8";
      when  650 => r := x"3ebf78313f9c8cf6";
      when  651 => r := x"3ebf3db33f9c750a";
      when  652 => r := x"3ebf03503f9c5d26";
      when  653 => r := x"3ebec9083f9c4549";
      when  654 => r := x"3ebe8eda3f9c2d74";
      when  655 => r := x"3ebe54c73f9c15a6";
      when  656 => r := x"3ebe1ace3f9bfddf";
      when  657 => r := x"3ebde0f03f9be61f";
      when  658 => r := x"3ebda72c3f9bce66";
      when  659 => r := x"3ebd6d833f9bb6b5";
      when  660 => r := x"3ebd33f43f9b9f0b";
      when  661 => r := x"3ebcfa7f3f9b8768";
      when  662 => r := x"3ebcc1243f9b6fcc";
      when  663 => r := x"3ebc87e43f9b5838";
      when  664 => r := x"3ebc4ebd3f9b40aa";
      when  665 => r := x"3ebc15b03f9b2924";
      when  666 => r := x"3ebbdcbe3f9b11a5";
      when  667 => r := x"3ebba3e53f9afa2d";
      when  668 => r := x"3ebb6b263f9ae2bc";
      when  669 => r := x"3ebb32803f9acb52";
      when  670 => r := x"3ebaf9f53f9ab3ef";
      when  671 => r := x"3ebac1823f9a9c94";
      when  672 => r := x"3eba892a3f9a853f";
      when  673 => r := x"3eba50eb3f9a6df1";
      when  674 => r := x"3eba18c53f9a56ab";
      when  675 => r := x"3eb9e0b93f9a3f6b";
      when  676 => r := x"3eb9a8c63f9a2833";
      when  677 => r := x"3eb970ec3f9a1101";
      when  678 => r := x"3eb9392c3f99f9d6";
      when  679 => r := x"3eb901843f99e2b3";
      when  680 => r := x"3eb8c9f63f99cb96";
      when  681 => r := x"3eb892813f99b480";
      when  682 => r := x"3eb85b243f999d71";
      when  683 => r := x"3eb823e13f998669";
      when  684 => r := x"3eb7ecb63f996f68";
      when  685 => r := x"3eb7b5a43f99586e";
      when  686 => r := x"3eb77eab3f99417b";
      when  687 => r := x"3eb747cb3f992a8f";
      when  688 => r := x"3eb711033f9913a9";
      when  689 => r := x"3eb6da533f98fcca";
      when  690 => r := x"3eb6a3bc3f98e5f2";
      when  691 => r := x"3eb66d3e3f98cf21";
      when  692 => r := x"3eb636d83f98b857";
      when  693 => r := x"3eb6008a3f98a194";
      when  694 => r := x"3eb5ca553f988ad7";
      when  695 => r := x"3eb594373f987421";
      when  696 => r := x"3eb55e323f985d72";
      when  697 => r := x"3eb528453f9846ca";
      when  698 => r := x"3eb4f2703f983028";
      when  699 => r := x"3eb4bcb33f98198d";
      when  700 => r := x"3eb4870e3f9802f9";
      when  701 => r := x"3eb451813f97ec6b";
      when  702 => r := x"3eb41c0c3f97d5e4";
      when  703 => r := x"3eb3e6ae3f97bf64";
      when  704 => r := x"3eb3b1683f97a8eb";
      when  705 => r := x"3eb37c3a3f979278";
      when  706 => r := x"3eb347233f977c0c";
      when  707 => r := x"3eb312243f9765a6";
      when  708 => r := x"3eb2dd3c3f974f47";
      when  709 => r := x"3eb2a86c3f9738ef";
      when  710 => r := x"3eb273b33f97229d";
      when  711 => r := x"3eb23f123f970c52";
      when  712 => r := x"3eb20a873f96f60d";
      when  713 => r := x"3eb1d6143f96dfcf";
      when  714 => r := x"3eb1a1b83f96c998";
      when  715 => r := x"3eb16d743f96b367";
      when  716 => r := x"3eb139463f969d3c";
      when  717 => r := x"3eb1052f3f968718";
      when  718 => r := x"3eb0d12f3f9670fb";
      when  719 => r := x"3eb09d473f965ae4";
      when  720 => r := x"3eb069753f9644d4";
      when  721 => r := x"3eb035b93f962eca";
      when  722 => r := x"3eb002153f9618c6";
      when  723 => r := x"3eafce873f9602c9";
      when  724 => r := x"3eaf9b103f95ecd3";
      when  725 => r := x"3eaf67af3f95d6e2";
      when  726 => r := x"3eaf34653f95c0f9";
      when  727 => r := x"3eaf01323f95ab15";
      when  728 => r := x"3eaece153f959538";
      when  729 => r := x"3eae9b0e3f957f62";
      when  730 => r := x"3eae681d3f956992";
      when  731 => r := x"3eae35433f9553c8";
      when  732 => r := x"3eae027f3f953e04";
      when  733 => r := x"3eadcfd23f952847";
      when  734 => r := x"3ead9d3a3f951290";
      when  735 => r := x"3ead6ab93f94fce0";
      when  736 => r := x"3ead384d3f94e736";
      when  737 => r := x"3ead05f83f94d192";
      when  738 => r := x"3eacd3b83f94bbf4";
      when  739 => r := x"3eaca18e3f94a65d";
      when  740 => r := x"3eac6f7a3f9490cc";
      when  741 => r := x"3eac3d7c3f947b41";
      when  742 => r := x"3eac0b943f9465bc";
      when  743 => r := x"3eabd9c13f94503e";
      when  744 => r := x"3eaba8043f943ac6";
      when  745 => r := x"3eab765d3f942554";
      when  746 => r := x"3eab44cb3f940fe8";
      when  747 => r := x"3eab134e3f93fa83";
      when  748 => r := x"3eaae1e73f93e523";
      when  749 => r := x"3eaab0963f93cfca";
      when  750 => r := x"3eaa7f593f93ba77";
      when  751 => r := x"3eaa4e323f93a52a";
      when  752 => r := x"3eaa1d203f938fe4";
      when  753 => r := x"3ea9ec243f937aa3";
      when  754 => r := x"3ea9bb3c3f936569";
      when  755 => r := x"3ea98a6a3f935034";
      when  756 => r := x"3ea959ad3f933b06";
      when  757 => r := x"3ea929053f9325de";
      when  758 => r := x"3ea8f8713f9310bc";
      when  759 => r := x"3ea8c7f33f92fba0";
      when  760 => r := x"3ea897893f92e68a";
      when  761 => r := x"3ea867353f92d17a";
      when  762 => r := x"3ea836f53f92bc70";
      when  763 => r := x"3ea806c93f92a76c";
      when  764 => r := x"3ea7d6b33f92926e";
      when  765 => r := x"3ea7a6b13f927d77";
      when  766 => r := x"3ea776c43f926885";
      when  767 => r := x"3ea746eb3f925399";
      when  768 => r := x"3ea717263f923eb3";
      when  769 => r := x"3ea6e7773f9229d3";
      when  770 => r := x"3ea6b7db3f9214f9";
      when  771 => r := x"3ea688543f920025";
      when  772 => r := x"3ea658e13f91eb57";
      when  773 => r := x"3ea629833f91d68f";
      when  774 => r := x"3ea5fa393f91c1cd";
      when  775 => r := x"3ea5cb023f91ad10";
      when  776 => r := x"3ea59be03f91985a";
      when  777 => r := x"3ea56cd33f9183a9";
      when  778 => r := x"3ea53dd93f916eff";
      when  779 => r := x"3ea50ef33f915a5a";
      when  780 => r := x"3ea4e0213f9145bb";
      when  781 => r := x"3ea4b1633f913122";
      when  782 => r := x"3ea482b93f911c8f";
      when  783 => r := x"3ea454233f910801";
      when  784 => r := x"3ea425a03f90f37a";
      when  785 => r := x"3ea3f7313f90def8";
      when  786 => r := x"3ea3c8d63f90ca7c";
      when  787 => r := x"3ea39a8f3f90b605";
      when  788 => r := x"3ea36c5b3f90a195";
      when  789 => r := x"3ea33e3b3f908d2a";
      when  790 => r := x"3ea3102e3f9078c5";
      when  791 => r := x"3ea2e2353f906466";
      when  792 => r := x"3ea2b44f3f90500d";
      when  793 => r := x"3ea2867c3f903bb9";
      when  794 => r := x"3ea258bd3f90276b";
      when  795 => r := x"3ea22b113f901323";
      when  796 => r := x"3ea1fd793f8ffee1";
      when  797 => r := x"3ea1cff33f8feaa4";
      when  798 => r := x"3ea1a2813f8fd66d";
      when  799 => r := x"3ea175223f8fc23b";
      when  800 => r := x"3ea147d63f8fae0f";
      when  801 => r := x"3ea11a9e3f8f99e9";
      when  802 => r := x"3ea0ed783f8f85c9";
      when  803 => r := x"3ea0c0653f8f71ae";
      when  804 => r := x"3ea093653f8f5d99";
      when  805 => r := x"3ea066783f8f4989";
      when  806 => r := x"3ea0399d3f8f357f";
      when  807 => r := x"3ea00cd63f8f217a";
      when  808 => r := x"3e9fe0213f8f0d7c";
      when  809 => r := x"3e9fb37f3f8ef982";
      when  810 => r := x"3e9f86f03f8ee58f";
      when  811 => r := x"3e9f5a733f8ed1a1";
      when  812 => r := x"3e9f2e093f8ebdb8";
      when  813 => r := x"3e9f01b23f8ea9d5";
      when  814 => r := x"3e9ed56d3f8e95f8";
      when  815 => r := x"3e9ea93b3f8e8220";
      when  816 => r := x"3e9e7d1a3f8e6e4d";
      when  817 => r := x"3e9e510d3f8e5a81";
      when  818 => r := x"3e9e25123f8e46b9";
      when  819 => r := x"3e9df9293f8e32f7";
      when  820 => r := x"3e9dcd523f8e1f3b";
      when  821 => r := x"3e9da18d3f8e0b84";
      when  822 => r := x"3e9d75db3f8df7d2";
      when  823 => r := x"3e9d4a3b3f8de426";
      when  824 => r := x"3e9d1ead3f8dd080";
      when  825 => r := x"3e9cf3313f8dbcdf";
      when  826 => r := x"3e9cc7c73f8da943";
      when  827 => r := x"3e9c9c6f3f8d95ad";
      when  828 => r := x"3e9c712a3f8d821c";
      when  829 => r := x"3e9c45f63f8d6e91";
      when  830 => r := x"3e9c1ad43f8d5b0b";
      when  831 => r := x"3e9befc33f8d478a";
      when  832 => r := x"3e9bc4c53f8d340f";
      when  833 => r := x"3e9b99d83f8d2099";
      when  834 => r := x"3e9b6efd3f8d0d28";
      when  835 => r := x"3e9b44343f8cf9bd";
      when  836 => r := x"3e9b197d3f8ce657";
      when  837 => r := x"3e9aeed73f8cd2f7";
      when  838 => r := x"3e9ac4423f8cbf9b";
      when  839 => r := x"3e9a99bf3f8cac45";
      when  840 => r := x"3e9a6f4e3f8c98f5";
      when  841 => r := x"3e9a44ee3f8c85aa";
      when  842 => r := x"3e9a1aa03f8c7264";
      when  843 => r := x"3e99f0633f8c5f23";
      when  844 => r := x"3e99c6373f8c4be8";
      when  845 => r := x"3e999c1d3f8c38b1";
      when  846 => r := x"3e9972143f8c2581";
      when  847 => r := x"3e99481c3f8c1255";
      when  848 => r := x"3e991e353f8bff2e";
      when  849 => r := x"3e98f4603f8bec0d";
      when  850 => r := x"3e98ca9c3f8bd8f1";
      when  851 => r := x"3e98a0e83f8bc5db";
      when  852 => r := x"3e9877463f8bb2c9";
      when  853 => r := x"3e984db53f8b9fbd";
      when  854 => r := x"3e9824353f8b8cb6";
      when  855 => r := x"3e97fac63f8b79b4";
      when  856 => r := x"3e97d1683f8b66b7";
      when  857 => r := x"3e97a81a3f8b53bf";
      when  858 => r := x"3e977ede3f8b40cd";
      when  859 => r := x"3e9755b23f8b2de0";
      when  860 => r := x"3e972c973f8b1af8";
      when  861 => r := x"3e97038d3f8b0815";
      when  862 => r := x"3e96da933f8af537";
      when  863 => r := x"3e96b1ab3f8ae25e";
      when  864 => r := x"3e9688d23f8acf8a";
      when  865 => r := x"3e96600b3f8abcbc";
      when  866 => r := x"3e9637543f8aa9f2";
      when  867 => r := x"3e960ead3f8a972e";
      when  868 => r := x"3e95e6173f8a846f";
      when  869 => r := x"3e95bd923f8a71b4";
      when  870 => r := x"3e95951c3f8a5eff";
      when  871 => r := x"3e956cb83f8a4c4f";
      when  872 => r := x"3e9544633f8a39a4";
      when  873 => r := x"3e951c1f3f8a26fe";
      when  874 => r := x"3e94f3eb3f8a145d";
      when  875 => r := x"3e94cbc83f8a01c1";
      when  876 => r := x"3e94a3b43f89ef2a";
      when  877 => r := x"3e947bb13f89dc98";
      when  878 => r := x"3e9453be3f89ca0b";
      when  879 => r := x"3e942bdb3f89b783";
      when  880 => r := x"3e9404093f89a500";
      when  881 => r := x"3e93dc463f899282";
      when  882 => r := x"3e93b4933f898009";
      when  883 => r := x"3e938cf03f896d95";
      when  884 => r := x"3e93655e3f895b26";
      when  885 => r := x"3e933ddb3f8948bc";
      when  886 => r := x"3e9316683f893656";
      when  887 => r := x"3e92ef043f8923f6";
      when  888 => r := x"3e92c7b13f89119b";
      when  889 => r := x"3e92a06d3f88ff44";
      when  890 => r := x"3e92793a3f88ecf2";
      when  891 => r := x"3e9252153f88daa6";
      when  892 => r := x"3e922b013f88c85e";
      when  893 => r := x"3e9203fc3f88b61b";
      when  894 => r := x"3e91dd073f88a3dd";
      when  895 => r := x"3e91b6213f8891a4";
      when  896 => r := x"3e918f4b3f887f6f";
      when  897 => r := x"3e9168853f886d40";
      when  898 => r := x"3e9141ce3f885b15";
      when  899 => r := x"3e911b263f8848ef";
      when  900 => r := x"3e90f48e3f8836cf";
      when  901 => r := x"3e90ce053f8824b2";
      when  902 => r := x"3e90a78c3f88129b";
      when  903 => r := x"3e9081223f880088";
      when  904 => r := x"3e905ac73f87ee7b";
      when  905 => r := x"3e90347b3f87dc72";
      when  906 => r := x"3e900e3f3f87ca6e";
      when  907 => r := x"3e8fe8123f87b86e";
      when  908 => r := x"3e8fc1f43f87a674";
      when  909 => r := x"3e8f9be53f87947e";
      when  910 => r := x"3e8f75e53f87828d";
      when  911 => r := x"3e8f4ff53f8770a0";
      when  912 => r := x"3e8f2a133f875eb9";
      when  913 => r := x"3e8f04413f874cd6";
      when  914 => r := x"3e8ede7d3f873af8";
      when  915 => r := x"3e8eb8c83f87291e";
      when  916 => r := x"3e8e93233f871749";
      when  917 => r := x"3e8e6d8c3f870579";
      when  918 => r := x"3e8e48043f86f3ae";
      when  919 => r := x"3e8e228b3f86e1e7";
      when  920 => r := x"3e8dfd203f86d025";
      when  921 => r := x"3e8dd7c53f86be68";
      when  922 => r := x"3e8db2783f86acaf";
      when  923 => r := x"3e8d8d3a3f869afb";
      when  924 => r := x"3e8d680a3f86894c";
      when  925 => r := x"3e8d42e93f8677a1";
      when  926 => r := x"3e8d1dd73f8665fb";
      when  927 => r := x"3e8cf8d43f86545a";
      when  928 => r := x"3e8cd3de3f8642bd";
      when  929 => r := x"3e8caef83f863125";
      when  930 => r := x"3e8c8a203f861f91";
      when  931 => r := x"3e8c65563f860e02";
      when  932 => r := x"3e8c409b3f85fc78";
      when  933 => r := x"3e8c1bee3f85eaf2";
      when  934 => r := x"3e8bf7503f85d971";
      when  935 => r := x"3e8bd2c03f85c7f4";
      when  936 => r := x"3e8bae3e3f85b67c";
      when  937 => r := x"3e8b89cb3f85a509";
      when  938 => r := x"3e8b65663f85939a";
      when  939 => r := x"3e8b410f3f85822f";
      when  940 => r := x"3e8b1cc63f8570ca";
      when  941 => r := x"3e8af88c3f855f68";
      when  942 => r := x"3e8ad45f3f854e0b";
      when  943 => r := x"3e8ab0413f853cb3";
      when  944 => r := x"3e8a8c313f852b5f";
      when  945 => r := x"3e8a682f3f851a10";
      when  946 => r := x"3e8a443a3f8508c5";
      when  947 => r := x"3e8a20543f84f77f";
      when  948 => r := x"3e89fc7c3f84e63d";
      when  949 => r := x"3e89d8b23f84d500";
      when  950 => r := x"3e89b4f63f84c3c7";
      when  951 => r := x"3e8991473f84b293";
      when  952 => r := x"3e896da73f84a163";
      when  953 => r := x"3e894a143f849037";
      when  954 => r := x"3e89268f3f847f10";
      when  955 => r := x"3e8903183f846dee";
      when  956 => r := x"3e88dfaf3f845ccf";
      when  957 => r := x"3e88bc533f844bb6";
      when  958 => r := x"3e8899053f843aa0";
      when  959 => r := x"3e8875c53f84298f";
      when  960 => r := x"3e8852933f841883";
      when  961 => r := x"3e882f6e3f84077b";
      when  962 => r := x"3e880c563f83f677";
      when  963 => r := x"3e87e94c3f83e578";
      when  964 => r := x"3e87c6503f83d47d";
      when  965 => r := x"3e87a3613f83c386";
      when  966 => r := x"3e8780803f83b294";
      when  967 => r := x"3e875dac3f83a1a6";
      when  968 => r := x"3e873ae53f8390bd";
      when  969 => r := x"3e87182c3f837fd7";
      when  970 => r := x"3e86f5803f836ef6";
      when  971 => r := x"3e86d2e23f835e1a";
      when  972 => r := x"3e86b0513f834d42";
      when  973 => r := x"3e868dcd3f833c6e";
      when  974 => r := x"3e866b573f832b9e";
      when  975 => r := x"3e8648ed3f831ad3";
      when  976 => r := x"3e8626913f830a0c";
      when  977 => r := x"3e8604423f82f949";
      when  978 => r := x"3e85e2003f82e88b";
      when  979 => r := x"3e85bfcc3f82d7d1";
      when  980 => r := x"3e859da43f82c71b";
      when  981 => r := x"3e857b8a3f82b669";
      when  982 => r := x"3e85597c3f82a5bc";
      when  983 => r := x"3e85377c3f829513";
      when  984 => r := x"3e8515893f82846e";
      when  985 => r := x"3e84f3a23f8273ce";
      when  986 => r := x"3e84d1c93f826331";
      when  987 => r := x"3e84affc3f825299";
      when  988 => r := x"3e848e3d3f824205";
      when  989 => r := x"3e846c8a3f823176";
      when  990 => r := x"3e844ae43f8220ea";
      when  991 => r := x"3e84294b3f821063";
      when  992 => r := x"3e8407bf3f81ffe0";
      when  993 => r := x"3e83e63f3f81ef61";
      when  994 => r := x"3e83c4cc3f81dee6";
      when  995 => r := x"3e83a3663f81ce70";
      when  996 => r := x"3e83820d3f81bdfd";
      when  997 => r := x"3e8360c03f81ad8f";
      when  998 => r := x"3e833f803f819d25";
      when  999 => r := x"3e831e4c3f818cbf";
      when 1000 => r := x"3e82fd253f817c5e";
      when 1001 => r := x"3e82dc0b3f816c00";
      when 1002 => r := x"3e82bafd3f815ba7";
      when 1003 => r := x"3e8299fc3f814b51";
      when 1004 => r := x"3e8279073f813b00";
      when 1005 => r := x"3e82581f3f812ab3";
      when 1006 => r := x"3e8237433f811a6a";
      when 1007 => r := x"3e8216743f810a25";
      when 1008 => r := x"3e81f5b13f80f9e5";
      when 1009 => r := x"3e81d4fa3f80e9a8";
      when 1010 => r := x"3e81b4503f80d96f";
      when 1011 => r := x"3e8193b23f80c93b";
      when 1012 => r := x"3e8173203f80b90a";
      when 1013 => r := x"3e81529b3f80a8de";
      when 1014 => r := x"3e8132213f8098b6";
      when 1015 => r := x"3e8111b43f808891";
      when 1016 => r := x"3e80f1543f807871";
      when 1017 => r := x"3e80d0ff3f806855";
      when 1018 => r := x"3e80b0b73f80583d";
      when 1019 => r := x"3e80907a3f804829";
      when 1020 => r := x"3e80704a3f803819";
      when 1021 => r := x"3e8050263f80280d";
      when 1022 => r := x"3e80300e3f801805";
      when 1023 => r := x"3e8010023f800801";
      when others => r := (others => '0');      -- 0 ~ 2047 まであるのであり得ない。
    end case;
    return r;
  end table;

  component fadd
    port(A : in  std_logic_vector(31 downto 0);
         B : in  std_logic_vector(31 downto 0);
         S : out std_logic_vector(31 downto 0));
  end component;

  component fmul
    port(A : in  std_logic_vector(31 downto 0);
         B : in  std_logic_vector(31 downto 0);
         S : out std_logic_vector(31 downto 0));
  end component; 
  
  constant nan   : std_logic_vector(31 downto 0) := x"7fffffff";
  constant zero  : std_logic_vector(31 downto 0) := x"00000000";
  constant nzero : std_logic_vector(31 downto 0) := x"80000000";
  constant inf   : std_logic_vector(31 downto 0) := x"7f800000";
  constant ninf  : std_logic_vector(31 downto 0) := x"ff800000";

  signal s1,s2,s3,s4,s5 : std_logic_vector(31 downto 0);

begin

  -- Component Instantiation
  fadd_connect : fadd port map(
    A => s3,
    B => s4,
    S => s5);

  fmul_connect : fmul port map(
    A => s1,
    B => s2,
    S => s3);

  do_finv : process(A, s1, s2, s3, s4, s5)
    variable org      : std_logic_vector(31 downto 0);
    variable result   : std_logic_vector(31 downto 0);
    variable fraction : std_logic_vector(31 downto 0);
    variable d        : std_logic_vector(7 downto 0);
    variable index    : std_logic_vector(10 downto 0);
    variable ab_unit  : std_logic_vector(63 downto 0);
    variable ka,kb,temp : std_logic_vector(31 downto 0);   --変更
  begin

    if is_metavalue(A) then
      S <= (others => 'X');
    else
      org := A;

      if (org(30 downto 23) = 255 and org(22 downto 0) /= 0) then
        result := nan;
      elsif org(31) = '0' and org(30 downto 23) = 0 then
        result := inf;
      elsif org(31) = '1' and org(30 downto 23) = 0 then
        result := ninf;
      elsif org = inf then
        result := zero;
      elsif org = ninf then
        result := nzero;
      else
        if org(22 downto 0) = 0 then
          result := org;
          if org(30 downto 23) >= 127 then
            d := org(30 downto 23) - 127;
            result(30 downto 23) := 127 - d;
          else
            d := 127 - org(30 downto 23);
            result(30 downto 23) := 127 + d;
          end if;
        else
          fraction := org;
          fraction(31) := '0';
          fraction(30 downto 23) := "01111111";
          index := fraction(22 downto 13);
          ab_unit := table(index);
          ka := ab_unit(63 downto 32);
          kb := ab_unit(31 downto 0);
          ka(31) := '1';

          s1 <= ka;
          s2 <= fraction;
          s4 <= kb;
          temp := s5;

          result(31) := org(31);
          if org(30 downto 23) >= 127 then
            d := org(30 downto 23) - 127;
            if d < 126 then
              result(30 downto 23) := 126 - d; -- 127 - d - 1
              result(22 downto 0)  := temp(22 downto 0);
            else
              result(30 downto 0) := "000" & x"0000000";
            end if;
          else
            d := 127 - org(30 downto 23);
            result(30 downto 23) := 126 + d; -- 127 + d - 1
            result(22 downto 0)  := temp(22 downto 0);
          end if;
        end if;
      end if;

      S <= result;

    end if;
  end process;
end blackbox;
